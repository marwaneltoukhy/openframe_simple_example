magic
tech sky130A
magscale 1 2
timestamp 1695807346
<< obsli1 >>
rect 1104 2159 102856 101745
<< obsm1 >>
rect 14 2128 102856 101776
<< metal2 >>
rect 63130 103200 63186 104000
rect 18 0 74 800
rect 81162 0 81218 800
<< obsm2 >>
rect 20 103144 63074 103306
rect 63242 103144 99986 103306
rect 20 856 99986 103144
rect 130 800 81106 856
rect 81274 800 99986 856
<< metal3 >>
rect 0 85008 800 85128
rect 103200 61208 104000 61328
<< obsm3 >>
rect 800 85208 103200 101761
rect 880 84928 103200 85208
rect 800 61408 103200 84928
rect 800 61128 103120 61408
rect 800 2143 103200 61128
<< metal4 >>
rect 4208 2128 4528 101776
rect 19568 2128 19888 101776
rect 34928 2128 35248 101776
rect 50288 2128 50608 101776
rect 65648 2128 65968 101776
rect 81008 2128 81328 101776
rect 96368 2128 96688 101776
<< labels >>
rlabel metal3 s 0 85008 800 85128 6 a
port 1 nsew signal input
rlabel metal2 s 18 0 74 800 6 b
port 2 nsew signal input
rlabel metal3 s 103200 61208 104000 61328 6 clk
port 3 nsew signal input
rlabel metal2 s 63130 103200 63186 104000 6 out
port 4 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 rst
port 5 nsew signal input
rlabel metal4 s 4208 2128 4528 101776 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 101776 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 101776 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 101776 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 101776 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 101776 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 101776 6 vssd1
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 104000 104000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2773016
string GDS_FILE /home/marwan/openframe_simple_example/openlane/simple_design/runs/23_09_27_12_34/results/signoff/simple_design.magic.gds
string GDS_START 58204
<< end >>

