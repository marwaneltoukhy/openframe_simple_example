magic
tech sky130A
magscale 1 2
timestamp 1694959044
<< obsli1 >>
rect 8004 8143 625324 944945
<< obsm1 >>
rect 2774 2660 629266 950020
<< metal2 >>
rect 27498 953270 27558 953590
rect 29498 953270 29558 953590
rect 34360 953270 34416 953750
rect 34912 953270 34968 953750
rect 35556 953270 35612 953750
rect 36200 953270 36256 953750
rect 38040 953270 38096 953750
rect 38592 953270 38648 953750
rect 39236 953270 39292 953750
rect 39880 953270 39936 953750
rect 42364 953270 42420 953750
rect 42916 953270 42972 953750
rect 43560 953270 43616 953750
rect 44204 953270 44260 953750
rect 44756 953270 44812 953750
rect 45400 953270 45456 953750
rect 46596 953270 46652 953750
rect 47240 953270 47296 953750
rect 49080 953270 49136 953750
rect 78698 953270 78758 953590
rect 80698 953270 80758 953590
rect 85760 953270 85816 953750
rect 86312 953270 86368 953750
rect 86956 953270 87012 953750
rect 87600 953270 87656 953750
rect 89440 953270 89496 953750
rect 89992 953270 90048 953750
rect 90636 953270 90692 953750
rect 91280 953270 91336 953750
rect 93764 953270 93820 953750
rect 94316 953270 94372 953750
rect 94960 953270 95016 953750
rect 95604 953270 95660 953750
rect 96156 953270 96212 953750
rect 96800 953270 96856 953750
rect 97996 953270 98052 953750
rect 98640 953270 98696 953750
rect 100480 953270 100536 953750
rect 129898 953270 129958 953590
rect 131898 953270 131958 953590
rect 137160 953270 137216 953750
rect 137712 953270 137768 953750
rect 138356 953270 138412 953750
rect 139000 953270 139056 953750
rect 140840 953270 140896 953750
rect 141392 953270 141448 953750
rect 142036 953270 142092 953750
rect 142680 953270 142736 953750
rect 145164 953270 145220 953750
rect 145716 953270 145772 953750
rect 146360 953270 146416 953750
rect 147004 953270 147060 953750
rect 147556 953270 147612 953750
rect 148200 953270 148256 953750
rect 149396 953270 149452 953750
rect 150040 953270 150096 953750
rect 151880 953270 151936 953750
rect 181098 953270 181158 953590
rect 183098 953270 183158 953590
rect 188560 953270 188616 953750
rect 189112 953270 189168 953750
rect 189756 953270 189812 953750
rect 190400 953270 190456 953750
rect 192240 953270 192296 953750
rect 192792 953270 192848 953750
rect 193436 953270 193492 953750
rect 194080 953270 194136 953750
rect 196564 953270 196620 953750
rect 197116 953270 197172 953750
rect 197760 953270 197816 953750
rect 198404 953270 198460 953750
rect 198956 953270 199012 953750
rect 199600 953270 199656 953750
rect 200796 953270 200852 953750
rect 201440 953270 201496 953750
rect 203280 953270 203336 953750
rect 232298 953270 232358 953590
rect 234298 953270 234358 953590
rect 240160 953270 240216 953750
rect 240712 953270 240768 953750
rect 241356 953270 241412 953750
rect 242000 953270 242056 953750
rect 243840 953270 243896 953750
rect 244392 953270 244448 953750
rect 245036 953270 245092 953750
rect 245680 953270 245736 953750
rect 248164 953270 248220 953750
rect 248716 953270 248772 953750
rect 249360 953270 249416 953750
rect 250004 953270 250060 953750
rect 250556 953270 250612 953750
rect 251200 953270 251256 953750
rect 252396 953270 252452 953750
rect 253040 953270 253096 953750
rect 254880 953270 254936 953750
rect 336698 953270 336758 953590
rect 338698 953270 338758 953590
rect 341960 953270 342016 953750
rect 342512 953270 342568 953750
rect 343156 953270 343212 953750
rect 343800 953270 343856 953750
rect 345640 953270 345696 953750
rect 346192 953270 346248 953750
rect 346836 953270 346892 953750
rect 347480 953270 347536 953750
rect 349964 953270 350020 953750
rect 350516 953270 350572 953750
rect 351160 953270 351216 953750
rect 351804 953270 351860 953750
rect 352356 953270 352412 953750
rect 353000 953270 353056 953750
rect 354196 953270 354252 953750
rect 354840 953270 354896 953750
rect 356680 953270 356736 953750
rect 425698 953270 425758 953590
rect 427698 953270 427758 953590
rect 430960 953270 431016 953750
rect 431512 953270 431568 953750
rect 432156 953270 432212 953750
rect 432800 953270 432856 953750
rect 434640 953270 434696 953750
rect 435192 953270 435248 953750
rect 435836 953270 435892 953750
rect 436480 953270 436536 953750
rect 438964 953270 439020 953750
rect 439516 953270 439572 953750
rect 440160 953270 440216 953750
rect 440804 953270 440860 953750
rect 441356 953270 441412 953750
rect 442000 953270 442056 953750
rect 443196 953270 443252 953750
rect 443840 953270 443896 953750
rect 445680 953270 445736 953750
rect 476898 953270 476958 953590
rect 478898 953270 478958 953590
rect 482360 953270 482416 953750
rect 482912 953270 482968 953750
rect 483556 953270 483612 953750
rect 484200 953270 484256 953750
rect 486040 953270 486096 953750
rect 486592 953270 486648 953750
rect 487236 953270 487292 953750
rect 487880 953270 487936 953750
rect 490364 953270 490420 953750
rect 490916 953270 490972 953750
rect 491560 953270 491616 953750
rect 492204 953270 492260 953750
rect 492756 953270 492812 953750
rect 493400 953270 493456 953750
rect 494596 953270 494652 953750
rect 495240 953270 495296 953750
rect 497080 953270 497136 953750
rect 576298 953270 576358 953590
rect 578298 953270 578358 953590
rect 584160 953270 584216 953750
rect 584712 953270 584768 953750
rect 585356 953270 585412 953750
rect 586000 953270 586056 953750
rect 587840 953270 587896 953750
rect 588392 953270 588448 953750
rect 589036 953270 589092 953750
rect 589680 953270 589736 953750
rect 592164 953270 592220 953750
rect 592716 953270 592772 953750
rect 593360 953270 593416 953750
rect 594004 953270 594060 953750
rect 594556 953270 594612 953750
rect 595200 953270 595256 953750
rect 596396 953270 596452 953750
rect 597040 953270 597096 953750
rect 598880 953270 598936 953750
rect 99571 -90 99637 56
rect 110164 -116 110220 56
rect 145190 -424 145246 56
rect 147030 -424 147086 56
rect 147674 -424 147730 56
rect 148870 -424 148926 56
rect 149514 -424 149570 56
rect 150066 -424 150122 56
rect 150710 -424 150766 56
rect 151354 -424 151410 56
rect 151906 -424 151962 56
rect 154390 -424 154446 56
rect 155034 -424 155090 56
rect 155678 -424 155734 56
rect 156230 -424 156286 56
rect 158070 -424 158126 56
rect 158714 -424 158770 56
rect 159358 -424 159414 56
rect 159910 -424 159966 56
rect 160580 -260 160632 56
rect 163791 -259 163843 57
rect 253790 -424 253846 56
rect 255630 -424 255686 56
rect 256274 -424 256330 56
rect 257470 -424 257526 56
rect 258114 -424 258170 56
rect 258666 -424 258722 56
rect 259310 -424 259366 56
rect 259954 -424 260010 56
rect 260506 -424 260562 56
rect 262990 -424 263046 56
rect 263634 -424 263690 56
rect 264278 -424 264334 56
rect 264830 -424 264886 56
rect 266670 -424 266726 56
rect 267314 -424 267370 56
rect 267958 -424 268014 56
rect 268510 -424 268566 56
rect 269180 -260 269232 56
rect 273360 -260 273412 56
rect 308590 -424 308646 56
rect 310430 -424 310486 56
rect 311074 -424 311130 56
rect 312270 -424 312326 56
rect 312914 -424 312970 56
rect 313466 -424 313522 56
rect 314110 -424 314166 56
rect 314754 -424 314810 56
rect 315306 -424 315362 56
rect 317790 -424 317846 56
rect 318434 -424 318490 56
rect 319078 -424 319134 56
rect 319630 -424 319686 56
rect 321470 -424 321526 56
rect 322114 -424 322170 56
rect 322758 -424 322814 56
rect 323310 -424 323366 56
rect 323980 -260 324032 56
rect 328165 -282 328217 34
rect 363390 -424 363446 56
rect 365230 -424 365286 56
rect 365874 -424 365930 56
rect 367070 -424 367126 56
rect 367714 -424 367770 56
rect 368266 -424 368322 56
rect 368910 -424 368966 56
rect 369554 -424 369610 56
rect 370106 -424 370162 56
rect 372590 -424 372646 56
rect 373234 -424 373290 56
rect 373878 -424 373934 56
rect 374430 -424 374486 56
rect 376270 -424 376326 56
rect 376914 -424 376970 56
rect 377558 -424 377614 56
rect 378110 -424 378166 56
rect 378780 -260 378832 56
rect 382978 -260 383030 56
rect 418190 -424 418246 56
rect 420030 -424 420086 56
rect 420674 -424 420730 56
rect 421870 -424 421926 56
rect 422514 -424 422570 56
rect 423066 -424 423122 56
rect 423710 -424 423766 56
rect 424354 -424 424410 56
rect 424906 -424 424962 56
rect 427390 -424 427446 56
rect 428034 -424 428090 56
rect 428678 -424 428734 56
rect 429230 -424 429286 56
rect 431070 -424 431126 56
rect 431714 -424 431770 56
rect 432358 -424 432414 56
rect 432910 -424 432966 56
rect 433580 -260 433632 56
rect 437778 -260 437830 56
rect 472990 -424 473046 56
rect 474830 -424 474886 56
rect 475474 -424 475530 56
rect 476670 -424 476726 56
rect 477314 -424 477370 56
rect 477866 -424 477922 56
rect 478510 -424 478566 56
rect 479154 -424 479210 56
rect 479706 -424 479762 56
rect 482190 -424 482246 56
rect 482834 -424 482890 56
rect 483478 -424 483534 56
rect 484030 -424 484086 56
rect 485870 -424 485926 56
rect 486514 -424 486570 56
rect 487158 -424 487214 56
rect 487710 -424 487766 56
rect 488380 -260 488432 56
rect 492635 -260 492687 56
rect 605082 -260 605134 56
rect 605306 -260 605358 56
rect 605530 -260 605582 56
rect 605754 -260 605806 56
rect 605978 -260 606030 56
rect 606202 -260 606254 56
rect 606426 -260 606478 56
rect 606650 -260 606702 56
rect 606874 -260 606926 56
rect 607098 -260 607150 56
rect 607322 -260 607374 56
rect 607546 -260 607598 56
rect 607770 -260 607822 56
rect 607994 -260 608046 56
rect 608218 -260 608270 56
rect 608442 -260 608494 56
rect 608666 -260 608718 56
rect 608890 -260 608942 56
rect 609114 -260 609166 56
rect 609338 -260 609390 56
rect 609562 -260 609614 56
rect 609786 -260 609838 56
rect 610010 -260 610062 56
rect 610234 -260 610286 56
rect 610458 -260 610510 56
rect 610682 -260 610734 56
rect 610906 -260 610958 56
rect 611130 -260 611182 56
rect 611354 -260 611406 56
rect 611578 -260 611630 56
rect 611802 -260 611854 56
rect 612026 -260 612078 56
<< obsm2 >>
rect 2778 953214 27442 953306
rect 27614 953214 29442 953306
rect 29614 953214 34304 953306
rect 34472 953214 34856 953306
rect 35024 953214 35500 953306
rect 35668 953214 36144 953306
rect 36312 953214 37984 953306
rect 38152 953214 38536 953306
rect 38704 953214 39180 953306
rect 39348 953214 39824 953306
rect 39992 953214 42308 953306
rect 42476 953214 42860 953306
rect 43028 953214 43504 953306
rect 43672 953214 44148 953306
rect 44316 953214 44700 953306
rect 44868 953214 45344 953306
rect 45512 953214 46540 953306
rect 46708 953214 47184 953306
rect 47352 953214 49024 953306
rect 49192 953214 78642 953306
rect 78814 953214 80642 953306
rect 80814 953214 85704 953306
rect 85872 953214 86256 953306
rect 86424 953214 86900 953306
rect 87068 953214 87544 953306
rect 87712 953214 89384 953306
rect 89552 953214 89936 953306
rect 90104 953214 90580 953306
rect 90748 953214 91224 953306
rect 91392 953214 93708 953306
rect 93876 953214 94260 953306
rect 94428 953214 94904 953306
rect 95072 953214 95548 953306
rect 95716 953214 96100 953306
rect 96268 953214 96744 953306
rect 96912 953214 97940 953306
rect 98108 953214 98584 953306
rect 98752 953214 100424 953306
rect 100592 953214 129842 953306
rect 130014 953214 131842 953306
rect 132014 953214 137104 953306
rect 137272 953214 137656 953306
rect 137824 953214 138300 953306
rect 138468 953214 138944 953306
rect 139112 953214 140784 953306
rect 140952 953214 141336 953306
rect 141504 953214 141980 953306
rect 142148 953214 142624 953306
rect 142792 953214 145108 953306
rect 145276 953214 145660 953306
rect 145828 953214 146304 953306
rect 146472 953214 146948 953306
rect 147116 953214 147500 953306
rect 147668 953214 148144 953306
rect 148312 953214 149340 953306
rect 149508 953214 149984 953306
rect 150152 953214 151824 953306
rect 151992 953214 181042 953306
rect 181214 953214 183042 953306
rect 183214 953214 188504 953306
rect 188672 953214 189056 953306
rect 189224 953214 189700 953306
rect 189868 953214 190344 953306
rect 190512 953214 192184 953306
rect 192352 953214 192736 953306
rect 192904 953214 193380 953306
rect 193548 953214 194024 953306
rect 194192 953214 196508 953306
rect 196676 953214 197060 953306
rect 197228 953214 197704 953306
rect 197872 953214 198348 953306
rect 198516 953214 198900 953306
rect 199068 953214 199544 953306
rect 199712 953214 200740 953306
rect 200908 953214 201384 953306
rect 201552 953214 203224 953306
rect 203392 953214 232242 953306
rect 232414 953214 234242 953306
rect 234414 953214 240104 953306
rect 240272 953214 240656 953306
rect 240824 953214 241300 953306
rect 241468 953214 241944 953306
rect 242112 953214 243784 953306
rect 243952 953214 244336 953306
rect 244504 953214 244980 953306
rect 245148 953214 245624 953306
rect 245792 953214 248108 953306
rect 248276 953214 248660 953306
rect 248828 953214 249304 953306
rect 249472 953214 249948 953306
rect 250116 953214 250500 953306
rect 250668 953214 251144 953306
rect 251312 953214 252340 953306
rect 252508 953214 252984 953306
rect 253152 953214 254824 953306
rect 254992 953214 336642 953306
rect 336814 953214 338642 953306
rect 338814 953214 341904 953306
rect 342072 953214 342456 953306
rect 342624 953214 343100 953306
rect 343268 953214 343744 953306
rect 343912 953214 345584 953306
rect 345752 953214 346136 953306
rect 346304 953214 346780 953306
rect 346948 953214 347424 953306
rect 347592 953214 349908 953306
rect 350076 953214 350460 953306
rect 350628 953214 351104 953306
rect 351272 953214 351748 953306
rect 351916 953214 352300 953306
rect 352468 953214 352944 953306
rect 353112 953214 354140 953306
rect 354308 953214 354784 953306
rect 354952 953214 356624 953306
rect 356792 953214 425642 953306
rect 425814 953214 427642 953306
rect 427814 953214 430904 953306
rect 431072 953214 431456 953306
rect 431624 953214 432100 953306
rect 432268 953214 432744 953306
rect 432912 953214 434584 953306
rect 434752 953214 435136 953306
rect 435304 953214 435780 953306
rect 435948 953214 436424 953306
rect 436592 953214 438908 953306
rect 439076 953214 439460 953306
rect 439628 953214 440104 953306
rect 440272 953214 440748 953306
rect 440916 953214 441300 953306
rect 441468 953214 441944 953306
rect 442112 953214 443140 953306
rect 443308 953214 443784 953306
rect 443952 953214 445624 953306
rect 445792 953214 476842 953306
rect 477014 953214 478842 953306
rect 479014 953214 482304 953306
rect 482472 953214 482856 953306
rect 483024 953214 483500 953306
rect 483668 953214 484144 953306
rect 484312 953214 485984 953306
rect 486152 953214 486536 953306
rect 486704 953214 487180 953306
rect 487348 953214 487824 953306
rect 487992 953214 490308 953306
rect 490476 953214 490860 953306
rect 491028 953214 491504 953306
rect 491672 953214 492148 953306
rect 492316 953214 492700 953306
rect 492868 953214 493344 953306
rect 493512 953214 494540 953306
rect 494708 953214 495184 953306
rect 495352 953214 497024 953306
rect 497192 953214 576242 953306
rect 576414 953214 578242 953306
rect 578414 953214 584104 953306
rect 584272 953214 584656 953306
rect 584824 953214 585300 953306
rect 585468 953214 585944 953306
rect 586112 953214 587784 953306
rect 587952 953214 588336 953306
rect 588504 953214 588980 953306
rect 589148 953214 589624 953306
rect 589792 953214 592108 953306
rect 592276 953214 592660 953306
rect 592828 953214 593304 953306
rect 593472 953214 593948 953306
rect 594116 953214 594500 953306
rect 594668 953214 595144 953306
rect 595312 953214 596340 953306
rect 596508 953214 596984 953306
rect 597152 953214 598824 953306
rect 598992 953214 629262 953306
rect 2778 113 629262 953214
rect 2778 112 163735 113
rect 2778 14 99515 112
rect 99693 14 110108 112
rect 110276 14 145134 112
rect 145302 14 146974 112
rect 147142 14 147618 112
rect 147786 14 148814 112
rect 148982 14 149458 112
rect 149626 14 150010 112
rect 150178 14 150654 112
rect 150822 14 151298 112
rect 151466 14 151850 112
rect 152018 14 154334 112
rect 154502 14 154978 112
rect 155146 14 155622 112
rect 155790 14 156174 112
rect 156342 14 158014 112
rect 158182 14 158658 112
rect 158826 14 159302 112
rect 159470 14 159854 112
rect 160022 14 160524 112
rect 160688 14 163735 112
rect 163899 112 629262 113
rect 163899 14 253734 112
rect 253902 14 255574 112
rect 255742 14 256218 112
rect 256386 14 257414 112
rect 257582 14 258058 112
rect 258226 14 258610 112
rect 258778 14 259254 112
rect 259422 14 259898 112
rect 260066 14 260450 112
rect 260618 14 262934 112
rect 263102 14 263578 112
rect 263746 14 264222 112
rect 264390 14 264774 112
rect 264942 14 266614 112
rect 266782 14 267258 112
rect 267426 14 267902 112
rect 268070 14 268454 112
rect 268622 14 269124 112
rect 269288 14 273304 112
rect 273468 14 308534 112
rect 308702 14 310374 112
rect 310542 14 311018 112
rect 311186 14 312214 112
rect 312382 14 312858 112
rect 313026 14 313410 112
rect 313578 14 314054 112
rect 314222 14 314698 112
rect 314866 14 315250 112
rect 315418 14 317734 112
rect 317902 14 318378 112
rect 318546 14 319022 112
rect 319190 14 319574 112
rect 319742 14 321414 112
rect 321582 14 322058 112
rect 322226 14 322702 112
rect 322870 14 323254 112
rect 323422 14 323924 112
rect 324088 90 363334 112
rect 324088 14 328109 90
rect 328273 14 363334 90
rect 363502 14 365174 112
rect 365342 14 365818 112
rect 365986 14 367014 112
rect 367182 14 367658 112
rect 367826 14 368210 112
rect 368378 14 368854 112
rect 369022 14 369498 112
rect 369666 14 370050 112
rect 370218 14 372534 112
rect 372702 14 373178 112
rect 373346 14 373822 112
rect 373990 14 374374 112
rect 374542 14 376214 112
rect 376382 14 376858 112
rect 377026 14 377502 112
rect 377670 14 378054 112
rect 378222 14 378724 112
rect 378888 14 382922 112
rect 383086 14 418134 112
rect 418302 14 419974 112
rect 420142 14 420618 112
rect 420786 14 421814 112
rect 421982 14 422458 112
rect 422626 14 423010 112
rect 423178 14 423654 112
rect 423822 14 424298 112
rect 424466 14 424850 112
rect 425018 14 427334 112
rect 427502 14 427978 112
rect 428146 14 428622 112
rect 428790 14 429174 112
rect 429342 14 431014 112
rect 431182 14 431658 112
rect 431826 14 432302 112
rect 432470 14 432854 112
rect 433022 14 433524 112
rect 433688 14 437722 112
rect 437886 14 472934 112
rect 473102 14 474774 112
rect 474942 14 475418 112
rect 475586 14 476614 112
rect 476782 14 477258 112
rect 477426 14 477810 112
rect 477978 14 478454 112
rect 478622 14 479098 112
rect 479266 14 479650 112
rect 479818 14 482134 112
rect 482302 14 482778 112
rect 482946 14 483422 112
rect 483590 14 483974 112
rect 484142 14 485814 112
rect 485982 14 486458 112
rect 486626 14 487102 112
rect 487270 14 487654 112
rect 487822 14 488324 112
rect 488488 14 492579 112
rect 492743 14 605026 112
rect 605190 14 605250 112
rect 605414 14 605474 112
rect 605638 14 605698 112
rect 605862 14 605922 112
rect 606086 14 606146 112
rect 606310 14 606370 112
rect 606534 14 606594 112
rect 606758 14 606818 112
rect 606982 14 607042 112
rect 607206 14 607266 112
rect 607430 14 607490 112
rect 607654 14 607714 112
rect 607878 14 607938 112
rect 608102 14 608162 112
rect 608326 14 608386 112
rect 608550 14 608610 112
rect 608774 14 608834 112
rect 608998 14 609058 112
rect 609222 14 609282 112
rect 609446 14 609506 112
rect 609670 14 609730 112
rect 609894 14 609954 112
rect 610118 14 610178 112
rect 610342 14 610402 112
rect 610566 14 610626 112
rect 610790 14 610850 112
rect 611014 14 611074 112
rect 611238 14 611298 112
rect 611462 14 611522 112
rect 611686 14 611746 112
rect 611910 14 611970 112
rect 612134 14 629262 112
<< metal3 >>
rect 633270 929007 633590 929069
rect -424 927073 56 927143
rect 633270 927005 633590 927067
rect -424 925233 56 925303
rect 633270 925103 633750 925173
rect -424 924589 56 924659
rect 633270 924551 633750 924621
rect 633270 923907 633750 923977
rect -424 923393 56 923463
rect 633270 923263 633750 923333
rect -424 922749 56 922819
rect -424 922197 56 922267
rect -424 921553 56 921623
rect 633270 921423 633750 921493
rect -424 920909 56 920979
rect 633270 920871 633750 920941
rect -424 920357 56 920427
rect 633270 920227 633750 920297
rect 633270 919583 633750 919653
rect -424 917873 56 917943
rect -424 917229 56 917299
rect 633270 917099 633750 917169
rect -424 916585 56 916655
rect 633270 916547 633750 916617
rect -424 916033 56 916103
rect 633270 915903 633750 915973
rect 633270 915259 633750 915329
rect 633270 914707 633750 914777
rect -424 914193 56 914263
rect 633270 914063 633750 914133
rect -424 913549 56 913619
rect -424 912905 56 912975
rect 633270 912867 633750 912937
rect -424 912353 56 912423
rect 633270 912223 633750 912293
rect 633270 910383 633750 910453
rect -264 906644 56 906704
rect -264 904644 56 904704
rect 633270 839007 633590 839069
rect 633270 837005 633590 837067
rect 633270 835903 633750 835973
rect 633270 835351 633750 835421
rect 633270 834707 633750 834777
rect 633270 834063 633750 834133
rect 633270 832223 633750 832293
rect 633270 831671 633750 831741
rect 633270 831027 633750 831097
rect 633270 830383 633750 830453
rect 633270 827899 633750 827969
rect 633270 827347 633750 827417
rect 633270 826703 633750 826773
rect 633270 826059 633750 826129
rect 633270 825507 633750 825577
rect 633270 824863 633750 824933
rect 633270 823667 633750 823737
rect 633270 823023 633750 823093
rect 633270 821183 633750 821253
rect -424 757273 56 757343
rect -424 755433 56 755503
rect -424 754789 56 754859
rect -424 753593 56 753663
rect -424 752949 56 753019
rect -424 752397 56 752467
rect -424 751753 56 751823
rect -424 751109 56 751179
rect -424 750557 56 750627
rect 633270 750007 633590 750069
rect -424 748073 56 748143
rect 633270 748005 633590 748067
rect -424 747429 56 747499
rect -424 746785 56 746855
rect 633270 746703 633750 746773
rect -424 746233 56 746303
rect 633270 746151 633750 746221
rect 633270 745507 633750 745577
rect 633270 744863 633750 744933
rect -424 744393 56 744463
rect -424 743749 56 743819
rect -424 743105 56 743175
rect 633270 743023 633750 743093
rect -424 742553 56 742623
rect 633270 742471 633750 742541
rect 633270 741827 633750 741897
rect 633270 741183 633750 741253
rect 633270 738699 633750 738769
rect 633270 738147 633750 738217
rect 633270 737503 633750 737573
rect 633270 736859 633750 736929
rect -264 736644 56 736704
rect 633270 736307 633750 736377
rect 633270 735663 633750 735733
rect -264 734644 56 734704
rect 633270 734467 633750 734537
rect 633270 733823 633750 733893
rect 633270 731983 633750 732053
rect -424 714073 56 714143
rect -424 712233 56 712303
rect -424 711589 56 711659
rect -424 710393 56 710463
rect -424 709749 56 709819
rect -424 709197 56 709267
rect -424 708553 56 708623
rect -424 707909 56 707979
rect -424 707357 56 707427
rect -424 704873 56 704943
rect 633270 705007 633590 705069
rect -424 704229 56 704299
rect -424 703585 56 703655
rect -424 703033 56 703103
rect 633270 703005 633590 703067
rect 633270 701703 633750 701773
rect -424 701193 56 701263
rect 633270 701151 633750 701221
rect -424 700549 56 700619
rect 633270 700507 633750 700577
rect -424 699905 56 699975
rect 633270 699863 633750 699933
rect -424 699353 56 699423
rect 633270 698023 633750 698093
rect 633270 697471 633750 697541
rect 633270 696827 633750 696897
rect 633270 696183 633750 696253
rect -264 693644 56 693704
rect 633270 693699 633750 693769
rect 633270 693147 633750 693217
rect 633270 692503 633750 692573
rect 633270 691859 633750 691929
rect -264 691644 56 691704
rect 633270 691307 633750 691377
rect 633270 690663 633750 690733
rect 633270 689467 633750 689537
rect 633270 688823 633750 688893
rect 633270 686983 633750 687053
rect -424 670873 56 670943
rect -424 669033 56 669103
rect -424 668389 56 668459
rect -424 667193 56 667263
rect -424 666549 56 666619
rect -424 665997 56 666067
rect -424 665353 56 665423
rect -424 664709 56 664779
rect -424 664157 56 664227
rect -424 661673 56 661743
rect -424 661029 56 661099
rect -424 660385 56 660455
rect 633270 660007 633590 660069
rect -424 659833 56 659903
rect -424 657993 56 658063
rect 633270 658005 633590 658067
rect -424 657349 56 657419
rect -424 656705 56 656775
rect 633270 656703 633750 656773
rect -424 656153 56 656223
rect 633270 656151 633750 656221
rect 633270 655507 633750 655577
rect 633270 654863 633750 654933
rect 633270 653023 633750 653093
rect 633270 652471 633750 652541
rect 633270 651827 633750 651897
rect 633270 651183 633750 651253
rect -264 650644 56 650704
rect -264 648644 56 648704
rect 633270 648699 633750 648769
rect 633270 648147 633750 648217
rect 633270 647503 633750 647573
rect 633270 646859 633750 646929
rect 633270 646307 633750 646377
rect 633270 645663 633750 645733
rect 633270 644467 633750 644537
rect 633270 643823 633750 643893
rect 633270 641983 633750 642053
rect -424 627673 56 627743
rect -424 625833 56 625903
rect -424 625189 56 625259
rect -424 623993 56 624063
rect -424 623349 56 623419
rect -424 622797 56 622867
rect -424 622153 56 622223
rect -424 621509 56 621579
rect -424 620957 56 621027
rect -424 618473 56 618543
rect -424 617829 56 617899
rect -424 617185 56 617255
rect -424 616633 56 616703
rect 633270 615007 633590 615069
rect -424 614793 56 614863
rect -424 614149 56 614219
rect -424 613505 56 613575
rect -424 612953 56 613023
rect 633270 613005 633590 613067
rect 633270 611503 633750 611573
rect 633270 610951 633750 611021
rect 633270 610307 633750 610377
rect 633270 609663 633750 609733
rect 633270 607823 633750 607893
rect -264 607644 56 607704
rect 633270 607271 633750 607341
rect 633270 606627 633750 606697
rect 633270 605983 633750 606053
rect -264 605644 56 605704
rect 633270 603499 633750 603569
rect 633270 602947 633750 603017
rect 633270 602303 633750 602373
rect 633270 601659 633750 601729
rect 633270 601107 633750 601177
rect 633270 600463 633750 600533
rect 633270 599267 633750 599337
rect 633270 598623 633750 598693
rect 633270 596783 633750 596853
rect -424 584473 56 584543
rect -424 582633 56 582703
rect -424 581989 56 582059
rect -424 580793 56 580863
rect -424 580149 56 580219
rect -424 579597 56 579667
rect -424 578953 56 579023
rect -424 578309 56 578379
rect -424 577757 56 577827
rect -424 575273 56 575343
rect -424 574629 56 574699
rect -424 573985 56 574055
rect -424 573433 56 573503
rect -424 571593 56 571663
rect -424 570949 56 571019
rect -424 570305 56 570375
rect 633270 570007 633590 570069
rect -424 569753 56 569823
rect 633270 568005 633590 568067
rect 633270 566503 633750 566573
rect 633270 565951 633750 566021
rect 633270 565307 633750 565377
rect -264 564644 56 564704
rect 633270 564663 633750 564733
rect 633270 562823 633750 562893
rect -264 562644 56 562704
rect 633270 562271 633750 562341
rect 633270 561627 633750 561697
rect 633270 560983 633750 561053
rect 633270 558499 633750 558569
rect 633270 557947 633750 558017
rect 633270 557303 633750 557373
rect 633270 556659 633750 556729
rect 633270 556107 633750 556177
rect 633270 555463 633750 555533
rect 633270 554267 633750 554337
rect 633270 553623 633750 553693
rect 633270 551783 633750 551853
rect -424 541273 56 541343
rect -424 539433 56 539503
rect -424 538789 56 538859
rect -424 537593 56 537663
rect -424 536949 56 537019
rect -424 536397 56 536467
rect -424 535753 56 535823
rect -424 535109 56 535179
rect -424 534557 56 534627
rect -424 532073 56 532143
rect -424 531429 56 531499
rect -424 530785 56 530855
rect -424 530233 56 530303
rect -424 528393 56 528463
rect -424 527749 56 527819
rect -424 527105 56 527175
rect -424 526553 56 526623
rect 633270 525007 633590 525069
rect 633270 523005 633590 523067
rect -264 521644 56 521704
rect 633270 521303 633750 521373
rect 633270 520751 633750 520821
rect 633270 520107 633750 520177
rect -264 519644 56 519704
rect 633270 519463 633750 519533
rect 633270 517623 633750 517693
rect 633270 517071 633750 517141
rect 633270 516427 633750 516497
rect 633270 515783 633750 515853
rect 633270 513299 633750 513369
rect 633270 512747 633750 512817
rect 633270 512103 633750 512173
rect 633270 511459 633750 511529
rect 633270 510907 633750 510977
rect 633270 510263 633750 510333
rect 633270 509067 633750 509137
rect 633270 508423 633750 508493
rect 633270 506583 633750 506653
rect -424 498073 56 498143
rect -424 496233 56 496303
rect -424 495589 56 495659
rect -424 494393 56 494463
rect -424 493749 56 493819
rect -424 493197 56 493267
rect -424 492553 56 492623
rect -424 491909 56 491979
rect -424 491357 56 491427
rect -424 488873 56 488943
rect -424 488229 56 488299
rect -424 487585 56 487655
rect -424 487033 56 487103
rect -424 485193 56 485263
rect -424 484549 56 484619
rect -424 483905 56 483975
rect -424 483353 56 483423
rect -264 478644 56 478704
rect -264 476644 56 476704
rect -424 370473 56 370543
rect -424 368633 56 368703
rect -424 367989 56 368059
rect -424 366793 56 366863
rect -424 366149 56 366219
rect -424 365597 56 365667
rect -424 364953 56 365023
rect -424 364309 56 364379
rect -424 363757 56 363827
rect -424 361273 56 361343
rect -424 360629 56 360699
rect -424 359985 56 360055
rect -424 359433 56 359503
rect -424 357593 56 357663
rect -424 356949 56 357019
rect -424 356305 56 356375
rect -424 355753 56 355823
rect -264 349644 56 349704
rect 633270 348007 633590 348069
rect -264 347644 56 347704
rect 633270 346005 633590 346067
rect 633270 344103 633750 344173
rect 633270 343551 633750 343621
rect 633270 342907 633750 342977
rect 633270 342263 633750 342333
rect 633270 340423 633750 340493
rect 633270 339871 633750 339941
rect 633270 339227 633750 339297
rect 633270 338583 633750 338653
rect 633270 336099 633750 336169
rect 633270 335547 633750 335617
rect 633270 334903 633750 334973
rect 633270 334259 633750 334329
rect 633270 333707 633750 333777
rect 633270 333063 633750 333133
rect 633270 331867 633750 331937
rect 633270 331223 633750 331293
rect 633270 329383 633750 329453
rect -424 327273 56 327343
rect -424 325433 56 325503
rect -424 324789 56 324859
rect -424 323593 56 323663
rect -424 322949 56 323019
rect -424 322397 56 322467
rect -424 321753 56 321823
rect -424 321109 56 321179
rect -424 320557 56 320627
rect -424 318073 56 318143
rect -424 317429 56 317499
rect -424 316785 56 316855
rect -424 316233 56 316303
rect -424 314393 56 314463
rect -424 313749 56 313819
rect -424 313105 56 313175
rect -424 312553 56 312623
rect -264 306644 56 306704
rect -264 304644 56 304704
rect 633270 303007 633590 303069
rect 633270 301005 633590 301067
rect 633270 298903 633750 298973
rect 633270 298351 633750 298421
rect 633270 297707 633750 297777
rect 633270 297063 633750 297133
rect 633270 295223 633750 295293
rect 633270 294671 633750 294741
rect 633270 294027 633750 294097
rect 633270 293383 633750 293453
rect 633270 290899 633750 290969
rect 633270 290347 633750 290417
rect 633270 289703 633750 289773
rect 633270 289059 633750 289129
rect 633270 288507 633750 288577
rect 633270 287863 633750 287933
rect 633270 286667 633750 286737
rect 633270 286023 633750 286093
rect -424 284073 56 284143
rect 633270 284183 633750 284253
rect -424 282233 56 282303
rect -424 281589 56 281659
rect -424 280393 56 280463
rect -424 279749 56 279819
rect -424 279197 56 279267
rect -424 278553 56 278623
rect -424 277909 56 277979
rect -424 277357 56 277427
rect -424 274873 56 274943
rect -424 274229 56 274299
rect -424 273585 56 273655
rect -424 273033 56 273103
rect -424 271193 56 271263
rect -424 270549 56 270619
rect -424 269905 56 269975
rect -424 269353 56 269423
rect -264 263644 56 263704
rect -264 261644 56 261704
rect 633270 258007 633590 258069
rect 633270 256005 633590 256067
rect 633270 253903 633750 253973
rect 633270 253351 633750 253421
rect 633270 252707 633750 252777
rect 633270 252063 633750 252133
rect 633270 250223 633750 250293
rect 633270 249671 633750 249741
rect 633270 249027 633750 249097
rect 633270 248383 633750 248453
rect 633270 245899 633750 245969
rect 633270 245347 633750 245417
rect 633270 244703 633750 244773
rect 633270 244059 633750 244129
rect 633270 243507 633750 243577
rect 633270 242863 633750 242933
rect 633270 241667 633750 241737
rect 633270 241023 633750 241093
rect -424 240873 56 240943
rect 633270 239183 633750 239253
rect -424 239033 56 239103
rect -424 238389 56 238459
rect -424 237193 56 237263
rect -424 236549 56 236619
rect -424 235997 56 236067
rect -424 235353 56 235423
rect -424 234709 56 234779
rect -424 234157 56 234227
rect -424 231673 56 231743
rect -424 231029 56 231099
rect -424 230385 56 230455
rect -424 229833 56 229903
rect -424 227993 56 228063
rect -424 227349 56 227419
rect -424 226705 56 226775
rect -424 226153 56 226223
rect -264 220644 56 220704
rect -264 218644 56 218704
rect 633270 213007 633590 213069
rect 633270 211005 633590 211067
rect 633270 208903 633750 208973
rect 633270 208351 633750 208421
rect 633270 207707 633750 207777
rect 633270 207063 633750 207133
rect 633270 205223 633750 205293
rect 633270 204671 633750 204741
rect 633270 204027 633750 204097
rect 633270 203383 633750 203453
rect 633270 200899 633750 200969
rect 633270 200347 633750 200417
rect 633270 199703 633750 199773
rect 633270 199059 633750 199129
rect 633270 198507 633750 198577
rect 633270 197863 633750 197933
rect -424 197672 56 197744
rect 633270 196667 633750 196737
rect 633270 196023 633750 196093
rect -424 195832 56 195904
rect -424 195188 56 195260
rect 633270 194183 633750 194253
rect -424 193992 56 194064
rect -424 193348 56 193420
rect -424 192796 56 192868
rect -424 192152 56 192224
rect -424 191508 56 191580
rect -424 190956 56 191028
rect -424 188472 56 188544
rect -424 187828 56 187900
rect -424 187184 56 187256
rect -424 186632 56 186704
rect -424 184792 56 184864
rect -424 184148 56 184220
rect -424 183504 56 183576
rect -424 182952 56 183024
rect -264 177644 56 177704
rect -264 175644 56 175704
rect 633270 168007 633590 168069
rect 633270 166005 633590 166067
rect 633270 163703 633750 163773
rect 633270 163151 633750 163221
rect 633270 162507 633750 162577
rect 633270 161863 633750 161933
rect 633270 160023 633750 160093
rect 633270 159471 633750 159541
rect 633270 158827 633750 158897
rect 633270 158183 633750 158253
rect 633270 155699 633750 155769
rect 633270 155147 633750 155217
rect -424 154472 56 154544
rect 633270 154503 633750 154573
rect 633270 153859 633750 153929
rect 633270 153307 633750 153377
rect -424 152632 56 152704
rect 633270 152663 633750 152733
rect -424 151988 56 152060
rect 633270 151467 633750 151537
rect -424 150792 56 150864
rect 633270 150823 633750 150893
rect -424 150148 56 150220
rect -424 149596 56 149668
rect -424 148952 56 149024
rect 633270 148983 633750 149053
rect -424 148308 56 148380
rect -424 147756 56 147828
rect -424 145272 56 145344
rect -424 144628 56 144700
rect -424 143984 56 144056
rect -424 143432 56 143504
rect -424 141592 56 141664
rect -424 140948 56 141020
rect -424 140304 56 140376
rect -424 139752 56 139824
rect -264 134644 56 134704
rect -264 132644 56 132704
rect 633270 123007 633590 123069
rect 633270 121005 633590 121067
rect 633270 118703 633750 118773
rect 633270 118151 633750 118221
rect 633270 117507 633750 117577
rect 633270 116863 633750 116933
rect 633270 115023 633750 115093
rect 633270 114471 633750 114541
rect 633270 113827 633750 113897
rect 633270 113183 633750 113253
rect 633270 110699 633750 110769
rect 633270 110147 633750 110217
rect 633270 109503 633750 109573
rect 633270 108859 633750 108929
rect 633270 108307 633750 108377
rect 633270 107663 633750 107733
rect 633270 106467 633750 106537
rect 633270 105823 633750 105893
rect 633270 103983 633750 104053
rect 633270 78007 633590 78069
rect 633270 76005 633590 76067
rect 633270 73503 633750 73573
rect 633270 72951 633750 73021
rect 633270 72307 633750 72377
rect 633270 71663 633750 71733
rect 633270 69823 633750 69893
rect 633270 69271 633750 69341
rect 633270 68627 633750 68697
rect 633270 67983 633750 68053
rect 633270 65499 633750 65569
rect 633270 64947 633750 65017
rect 633270 64303 633750 64373
rect 633270 63659 633750 63729
rect 633270 63107 633750 63177
rect 633270 62463 633750 62533
rect 633270 61267 633750 61337
rect 633270 60623 633750 60693
rect 633270 58783 633750 58853
rect -284 53595 56 53665
rect -284 53372 56 53442
rect -284 53147 56 53217
<< obsm3 >>
rect 0 929250 633326 944961
rect 0 929149 633328 929250
rect 0 928927 633190 929149
rect 633268 929114 633328 929149
rect 633206 929069 633328 929114
rect 0 927223 633326 928927
rect 136 927147 633326 927223
rect 136 926993 633190 927147
rect 0 926925 633190 926993
rect 0 925383 633326 926925
rect 136 925253 633326 925383
rect 136 925153 633190 925253
rect 0 925023 633190 925153
rect 0 924739 633326 925023
rect 136 924701 633326 924739
rect 136 924509 633190 924701
rect 0 924471 633190 924509
rect 0 924057 633326 924471
rect 0 923827 633190 924057
rect 0 923543 633326 923827
rect 136 923413 633326 923543
rect 136 923313 633190 923413
rect 0 923183 633190 923313
rect 0 922899 633326 923183
rect 136 922669 633326 922899
rect 0 922347 633326 922669
rect 136 922117 633326 922347
rect 0 921703 633326 922117
rect 136 921573 633326 921703
rect 136 921473 633190 921573
rect 0 921343 633190 921473
rect 0 921059 633326 921343
rect 136 921021 633326 921059
rect 136 920829 633190 921021
rect 0 920791 633190 920829
rect 0 920507 633326 920791
rect 136 920377 633326 920507
rect 136 920277 633190 920377
rect 0 920147 633190 920277
rect 0 919733 633326 920147
rect 0 919503 633190 919733
rect 0 918023 633326 919503
rect 136 917793 633326 918023
rect 0 917379 633326 917793
rect 136 917249 633326 917379
rect 136 917149 633190 917249
rect 0 917019 633190 917149
rect 0 917010 633326 917019
rect 0 916735 633328 917010
rect 136 916678 633328 916735
rect 136 916505 633190 916678
rect 0 916467 633190 916505
rect 0 916183 633326 916467
rect 136 916053 633326 916183
rect -2 915998 122 916033
rect -2 915953 58 915998
rect 136 915953 633190 916053
rect -2 915862 633190 915953
rect 0 915823 633190 915862
rect 0 915409 633326 915823
rect 0 915179 633190 915409
rect 0 914857 633326 915179
rect 0 914627 633190 914857
rect 0 914343 633326 914627
rect 136 914213 633326 914343
rect 136 914113 633190 914213
rect 0 913983 633190 914113
rect 0 913699 633326 913983
rect 136 913469 633326 913699
rect 0 913055 633326 913469
rect 136 913017 633326 913055
rect 136 912825 633190 913017
rect 0 912787 633190 912825
rect 0 912503 633326 912787
rect 136 912373 633326 912503
rect 136 912273 633190 912373
rect 0 912143 633190 912273
rect 0 910533 633326 912143
rect 0 910303 633190 910533
rect 0 906784 633326 910303
rect 136 906564 633326 906784
rect 0 904784 633326 906564
rect 136 904564 633326 904784
rect 0 880363 633326 904564
rect 0 865523 633571 880363
rect 0 839149 633326 865523
rect 0 838927 633190 839149
rect 0 837147 633326 838927
rect 0 836925 633190 837147
rect 0 836053 633326 836925
rect 0 835823 633190 836053
rect 0 835501 633326 835823
rect 0 835271 633190 835501
rect 0 834857 633326 835271
rect 0 834627 633190 834857
rect 0 834458 633326 834627
rect 0 834213 633328 834458
rect 0 833983 633190 834213
rect 633268 834186 633328 834213
rect 633206 834133 633328 834186
rect 0 832373 633326 833983
rect 0 832143 633190 832373
rect 0 831821 633326 832143
rect 0 831591 633190 831821
rect 0 831177 633326 831591
rect 0 830947 633190 831177
rect 0 830533 633326 830947
rect 0 830303 633190 830533
rect 0 828049 633326 830303
rect 0 827819 633190 828049
rect 0 827497 633326 827819
rect 0 827267 633190 827497
rect 0 826853 633326 827267
rect 0 826623 633190 826853
rect 0 826298 633326 826623
rect 0 826209 633328 826298
rect 0 825979 633190 826209
rect 633268 826162 633328 826209
rect 633206 826129 633328 826162
rect 0 825657 633326 825979
rect 0 825427 633190 825657
rect 0 825013 633326 825427
rect 0 824783 633190 825013
rect 0 823817 633326 824783
rect 0 823587 633190 823817
rect 0 823173 633326 823587
rect 0 822943 633190 823173
rect 633206 822974 633328 823023
rect 633268 822943 633328 822974
rect 0 822838 633328 822943
rect 0 821333 633326 822838
rect 0 821103 633190 821333
rect 0 757423 633326 821103
rect 136 757193 633326 757423
rect 0 755583 633326 757193
rect 136 755353 633326 755583
rect 0 754939 633326 755353
rect 136 754709 633326 754939
rect 0 753743 633326 754709
rect 136 753513 633326 753743
rect 0 753099 633326 753513
rect 136 752869 633326 753099
rect 0 752547 633326 752869
rect 136 752317 633326 752547
rect 0 751903 633326 752317
rect 136 751673 633326 751903
rect 0 751259 633326 751673
rect 136 751029 633326 751259
rect 0 750707 633326 751029
rect 136 750477 633326 750707
rect 0 750149 633326 750477
rect 0 749927 633190 750149
rect 0 748234 633326 749927
rect 0 748223 633328 748234
rect 136 748147 633328 748223
rect 136 747993 633190 748147
rect 633268 748098 633328 748147
rect 633206 748067 633328 748098
rect 0 747925 633190 747993
rect 0 747579 633326 747925
rect 136 747349 633326 747579
rect 0 746935 633326 747349
rect 136 746853 633326 746935
rect 136 746705 633190 746853
rect 0 746623 633190 746705
rect 0 746383 633326 746623
rect 136 746301 633326 746383
rect 136 746153 633190 746301
rect 0 746071 633190 746153
rect 0 745657 633326 746071
rect 0 745427 633190 745657
rect 0 745106 633326 745427
rect 0 745013 633328 745106
rect 0 744783 633190 745013
rect 633268 744970 633328 745013
rect 633206 744933 633328 744970
rect 0 744543 633326 744783
rect 136 744313 633326 744543
rect 0 743899 633326 744313
rect 136 743669 633326 743899
rect 0 743255 633326 743669
rect 136 743173 633326 743255
rect 136 743025 633190 743173
rect 0 742943 633190 743025
rect 0 742703 633326 742943
rect 136 742621 633326 742703
rect 136 742473 633190 742621
rect 0 742391 633190 742473
rect 0 741977 633326 742391
rect 0 741747 633190 741977
rect 0 741333 633326 741747
rect 0 741103 633190 741333
rect 0 738849 633326 741103
rect 0 738619 633190 738849
rect 0 738297 633326 738619
rect 0 738067 633190 738297
rect 633206 738110 633328 738147
rect 633268 738067 633328 738110
rect 0 737974 633328 738067
rect 0 737762 633326 737974
rect 0 737653 633328 737762
rect 0 737423 633190 737653
rect 633268 737626 633328 737653
rect 633206 737573 633328 737626
rect 0 737009 633326 737423
rect 0 736784 633190 737009
rect 136 736779 633190 736784
rect 136 736564 633326 736779
rect 0 736457 633326 736564
rect 0 736227 633190 736457
rect 0 735813 633326 736227
rect 0 735583 633190 735813
rect 0 734784 633326 735583
rect 136 734617 633326 734784
rect 136 734564 633190 734617
rect 0 734387 633190 734564
rect 0 733973 633326 734387
rect 0 733743 633190 733973
rect 0 732133 633326 733743
rect 0 731903 633190 732133
rect 0 714223 633326 731903
rect 136 713993 633326 714223
rect 0 712383 633326 713993
rect 136 712153 633326 712383
rect 0 711739 633326 712153
rect 136 711509 633326 711739
rect 0 710543 633326 711509
rect 136 710313 633326 710543
rect 0 709899 633326 710313
rect 136 709669 633326 709899
rect 0 709347 633326 709669
rect 136 709117 633326 709347
rect 0 708794 633326 709117
rect -2 708703 633326 708794
rect -2 708658 58 708703
rect -2 708623 122 708658
rect 136 708473 633326 708703
rect 0 708059 633326 708473
rect 136 707829 633326 708059
rect 0 707507 633326 707829
rect 136 707277 633326 707507
rect 0 705149 633326 707277
rect 0 705122 633190 705149
rect -2 705023 633190 705122
rect -2 704986 58 705023
rect -2 704943 122 704986
rect 136 704927 633190 705023
rect 136 704793 633326 704927
rect 0 704379 633326 704793
rect 136 704149 633326 704379
rect 0 703735 633326 704149
rect 136 703505 633326 703735
rect 0 703183 633326 703505
rect 136 703147 633326 703183
rect 136 702953 633190 703147
rect 0 702925 633190 702953
rect 0 701853 633326 702925
rect 0 701623 633190 701853
rect 0 701343 633326 701623
rect 136 701301 633326 701343
rect 136 701113 633190 701301
rect 0 701071 633190 701113
rect 0 700699 633326 701071
rect 136 700657 633326 700699
rect 136 700469 633190 700657
rect 0 700427 633190 700469
rect 0 700055 633326 700427
rect 136 700013 633326 700055
rect 136 699825 633190 700013
rect 0 699783 633190 699825
rect 0 699503 633326 699783
rect 136 699273 633326 699503
rect 0 698173 633326 699273
rect 0 697943 633190 698173
rect 633206 697990 633328 698023
rect 633268 697943 633328 697990
rect 0 697854 633328 697943
rect 0 697621 633326 697854
rect 0 697391 633190 697621
rect 0 696977 633326 697391
rect 0 696747 633190 696977
rect 0 696333 633326 696747
rect 0 696103 633190 696333
rect 0 693849 633326 696103
rect 0 693784 633190 693849
rect 136 693619 633190 693784
rect 136 693564 633326 693619
rect 0 693297 633326 693564
rect 0 693067 633190 693297
rect 0 692746 633326 693067
rect 0 692653 633328 692746
rect 0 692423 633190 692653
rect 633268 692610 633328 692653
rect 633206 692573 633328 692610
rect 0 692009 633326 692423
rect 0 691784 633190 692009
rect 136 691779 633190 691784
rect 136 691564 633326 691779
rect 0 691457 633326 691564
rect 0 691227 633190 691457
rect 0 690813 633326 691227
rect 0 690583 633190 690813
rect 0 689617 633326 690583
rect 0 689387 633190 689617
rect 0 688973 633326 689387
rect 0 688743 633190 688973
rect 0 687133 633326 688743
rect 0 686903 633190 687133
rect 0 671023 633326 686903
rect 136 670793 633326 671023
rect 0 669183 633326 670793
rect 136 668953 633326 669183
rect 0 668539 633326 668953
rect 136 668309 633326 668539
rect 0 667450 633326 668309
rect -2 667343 633326 667450
rect -2 667314 58 667343
rect -2 667263 122 667314
rect 136 667113 633326 667343
rect 0 666699 633326 667113
rect 136 666469 633326 666699
rect 0 666147 633326 666469
rect 136 665917 633326 666147
rect 0 665503 633326 665917
rect 136 665273 633326 665503
rect 0 664859 633326 665273
rect 136 664629 633326 664859
rect 0 664307 633326 664629
rect -2 664126 122 664157
rect -2 664077 58 664126
rect 136 664077 633326 664307
rect -2 663990 633326 664077
rect 0 661823 633326 663990
rect 136 661593 633326 661823
rect 0 661179 633326 661593
rect 136 660949 633326 661179
rect 0 660535 633326 660949
rect 136 660305 633326 660535
rect 0 660149 633326 660305
rect 0 659983 633190 660149
rect 136 659927 633190 659983
rect 136 659753 633326 659927
rect 0 658147 633326 659753
rect 0 658143 633190 658147
rect 136 657925 633190 658143
rect 136 657913 633326 657925
rect 0 657499 633326 657913
rect 136 657269 633326 657499
rect 0 656855 633326 657269
rect 136 656853 633326 656855
rect 136 656625 633190 656853
rect 0 656623 633190 656625
rect 0 656303 633326 656623
rect 136 656301 633326 656303
rect 136 656073 633190 656301
rect 0 656071 633190 656073
rect 0 655657 633326 656071
rect 0 655427 633190 655657
rect 0 655013 633326 655427
rect 0 654783 633190 655013
rect 0 653173 633326 654783
rect 0 652943 633190 653173
rect 0 652621 633326 652943
rect 0 652391 633190 652621
rect 0 651977 633326 652391
rect 0 651747 633190 651977
rect 0 651333 633326 651747
rect 0 651103 633190 651333
rect 0 650784 633326 651103
rect 136 650564 633326 650784
rect 0 648954 633326 650564
rect 0 648849 633328 648954
rect 0 648784 633190 648849
rect 633268 648818 633328 648849
rect 136 648619 633190 648784
rect 633206 648769 633328 648818
rect 136 648564 633326 648619
rect 0 648297 633326 648564
rect 0 648067 633190 648297
rect 0 647653 633326 648067
rect 0 647423 633190 647653
rect 0 647009 633326 647423
rect 0 646779 633190 647009
rect 0 646457 633326 646779
rect 0 646227 633190 646457
rect 0 645813 633326 646227
rect 0 645583 633190 645813
rect 633206 645630 633328 645663
rect 633268 645583 633328 645630
rect 0 645494 633328 645583
rect 0 644617 633326 645494
rect 0 644387 633190 644617
rect 0 643973 633326 644387
rect 0 643743 633190 643973
rect 0 642133 633326 643743
rect 0 641903 633190 642133
rect 0 627823 633326 641903
rect 136 627593 633326 627823
rect 0 625983 633326 627593
rect 136 625753 633326 625983
rect 0 625339 633326 625753
rect 136 625109 633326 625339
rect 0 624143 633326 625109
rect 136 623913 633326 624143
rect 0 623499 633326 623913
rect 136 623269 633326 623499
rect 0 622947 633326 623269
rect 136 622717 633326 622947
rect 0 622303 633326 622717
rect 136 622073 633326 622303
rect 0 621754 633326 622073
rect -2 621659 633326 621754
rect -2 621618 58 621659
rect -2 621579 122 621618
rect 136 621429 633326 621659
rect 0 621107 633326 621429
rect 136 620877 633326 621107
rect 0 618623 633326 620877
rect 136 618393 633326 618623
rect 0 617979 633326 618393
rect 136 617749 633326 617979
rect 0 617335 633326 617749
rect 136 617105 633326 617335
rect 0 616783 633326 617105
rect 136 616553 633326 616783
rect 0 615149 633326 616553
rect 0 614943 633190 615149
rect 136 614927 633190 614943
rect 136 614713 633326 614927
rect 0 614299 633326 614713
rect 136 614069 633326 614299
rect 0 613655 633326 614069
rect 136 613425 633326 613655
rect 0 613147 633326 613425
rect 0 613103 633190 613147
rect 136 612925 633190 613103
rect 136 612873 633326 612925
rect 0 611653 633326 612873
rect 0 611423 633190 611653
rect 0 611101 633326 611423
rect 0 610871 633190 611101
rect 0 610457 633326 610871
rect 0 610227 633190 610457
rect 633206 610270 633328 610307
rect 633268 610227 633328 610270
rect 0 610134 633328 610227
rect 0 609922 633326 610134
rect 0 609813 633328 609922
rect 0 609583 633190 609813
rect 633268 609786 633328 609813
rect 633206 609733 633328 609786
rect 0 607973 633326 609583
rect 0 607784 633190 607973
rect 136 607743 633190 607784
rect 136 607564 633326 607743
rect 0 607421 633326 607564
rect 0 607191 633190 607421
rect 0 606777 633326 607191
rect 0 606547 633190 606777
rect 0 606133 633326 606547
rect 0 605903 633190 606133
rect 0 605784 633326 605903
rect 136 605564 633326 605784
rect 0 603649 633326 605564
rect 0 603419 633190 603649
rect 0 603097 633326 603419
rect 0 602867 633190 603097
rect 0 602453 633326 602867
rect 0 602223 633190 602453
rect 0 601809 633326 602223
rect 0 601579 633190 601809
rect 0 601257 633326 601579
rect 0 601027 633190 601257
rect 0 600613 633326 601027
rect 0 600383 633190 600613
rect 0 599417 633326 600383
rect 0 599187 633190 599417
rect 0 598773 633326 599187
rect 0 598543 633190 598773
rect 0 596933 633326 598543
rect 0 596703 633190 596933
rect 0 584623 633326 596703
rect -2 584430 122 584473
rect -2 584393 58 584430
rect 136 584393 633326 584623
rect -2 584294 633326 584393
rect 0 582783 633326 584294
rect 136 582553 633326 582783
rect 0 582139 633326 582553
rect 136 581909 633326 582139
rect 0 580943 633326 581909
rect -2 580758 122 580793
rect -2 580713 58 580758
rect 136 580713 633326 580943
rect -2 580622 633326 580713
rect 0 580299 633326 580622
rect 136 580069 633326 580299
rect 0 579747 633326 580069
rect 136 579517 633326 579747
rect 0 579103 633326 579517
rect 136 578873 633326 579103
rect 0 578459 633326 578873
rect 136 578229 633326 578459
rect 0 577907 633326 578229
rect 136 577677 633326 577907
rect 0 575423 633326 577677
rect 136 575193 633326 575423
rect 0 574779 633326 575193
rect 136 574549 633326 574779
rect 0 574135 633326 574549
rect 136 573905 633326 574135
rect 0 573583 633326 573905
rect 136 573353 633326 573583
rect 0 571743 633326 573353
rect 136 571513 633326 571743
rect 0 571099 633326 571513
rect 136 570869 633326 571099
rect 0 570455 633326 570869
rect 136 570225 633326 570455
rect 0 570149 633326 570225
rect 0 569927 633190 570149
rect 0 569903 633326 569927
rect 136 569673 633326 569903
rect 0 568147 633326 569673
rect 0 567925 633190 568147
rect 633206 567974 633328 568005
rect 633268 567925 633328 567974
rect 0 567838 633328 567925
rect 0 566653 633326 567838
rect 0 566423 633190 566653
rect 0 566101 633326 566423
rect 0 565871 633190 566101
rect 0 565457 633326 565871
rect 0 565227 633190 565457
rect 0 564813 633326 565227
rect 0 564784 633190 564813
rect 136 564583 633190 564784
rect 136 564564 633326 564583
rect 0 562973 633326 564564
rect 0 562784 633190 562973
rect 136 562743 633190 562784
rect 136 562564 633326 562743
rect 0 562421 633326 562564
rect 0 562191 633190 562421
rect 0 561777 633326 562191
rect 0 561547 633190 561777
rect 0 561133 633326 561547
rect 0 560903 633190 561133
rect 0 558649 633326 560903
rect 0 558419 633190 558649
rect 0 558097 633326 558419
rect 0 557867 633190 558097
rect 0 557453 633326 557867
rect 0 557223 633190 557453
rect 0 556809 633326 557223
rect 0 556579 633190 556809
rect 0 556257 633326 556579
rect 0 556027 633190 556257
rect 0 555613 633326 556027
rect 0 555383 633190 555613
rect 0 554417 633326 555383
rect 0 554187 633190 554417
rect 0 553773 633326 554187
rect 0 553543 633190 553773
rect 0 551933 633326 553543
rect 0 551703 633190 551933
rect 0 541423 633326 551703
rect 136 541193 633326 541423
rect 0 539583 633326 541193
rect 136 539353 633326 539583
rect 0 538939 633326 539353
rect 136 538709 633326 538939
rect 0 537743 633326 538709
rect 136 537513 633326 537743
rect 0 537099 633326 537513
rect 136 536869 633326 537099
rect 0 536547 633326 536869
rect 136 536317 633326 536547
rect 0 535903 633326 536317
rect 136 535673 633326 535903
rect 0 535259 633326 535673
rect 136 535029 633326 535259
rect 0 534707 633326 535029
rect 136 534477 633326 534707
rect 0 532223 633326 534477
rect 136 531993 633326 532223
rect 0 531579 633326 531993
rect 136 531349 633326 531579
rect 0 530935 633326 531349
rect 136 530705 633326 530935
rect 0 530383 633326 530705
rect 136 530153 633326 530383
rect 0 528543 633326 530153
rect 136 528313 633326 528543
rect 0 527899 633326 528313
rect 136 527669 633326 527899
rect 0 527255 633326 527669
rect 136 527025 633326 527255
rect 0 526703 633326 527025
rect 136 526473 633326 526703
rect 0 525149 633326 526473
rect 0 524927 633190 525149
rect 0 523147 633326 524927
rect 0 522925 633190 523147
rect 0 521784 633326 522925
rect 136 521564 633326 521784
rect 0 521453 633326 521564
rect 0 521223 633190 521453
rect 0 520901 633326 521223
rect 0 520671 633190 520901
rect 0 520257 633326 520671
rect 0 520027 633190 520257
rect 0 519784 633326 520027
rect 136 519613 633326 519784
rect 136 519564 633190 519613
rect 0 519383 633190 519564
rect 0 517773 633326 519383
rect 0 517543 633190 517773
rect 0 517221 633326 517543
rect 0 516991 633190 517221
rect 0 516577 633326 516991
rect 0 516347 633190 516577
rect 0 515933 633326 516347
rect 0 515703 633190 515933
rect 633206 515750 633328 515783
rect 633268 515703 633328 515750
rect 0 515614 633328 515703
rect 0 513449 633326 515614
rect 0 513219 633190 513449
rect 0 512897 633326 513219
rect 0 512667 633190 512897
rect 0 512253 633326 512667
rect 0 512023 633190 512253
rect 0 511609 633326 512023
rect 0 511379 633190 511609
rect 0 511057 633326 511379
rect 0 510827 633190 511057
rect 0 510413 633326 510827
rect 0 510183 633190 510413
rect 0 509217 633326 510183
rect 0 508987 633190 509217
rect 0 508573 633326 508987
rect 0 508343 633190 508573
rect 0 506733 633326 508343
rect 0 506503 633190 506733
rect 0 498223 633326 506503
rect 136 497993 633326 498223
rect 0 496383 633326 497993
rect 136 496153 633326 496383
rect 0 495739 633326 496153
rect 136 495509 633326 495739
rect 0 494543 633326 495509
rect 136 494313 633326 494543
rect 0 493899 633326 494313
rect 136 493669 633326 493899
rect 0 493347 633326 493669
rect 136 493117 633326 493347
rect 0 492703 633326 493117
rect 136 492473 633326 492703
rect 0 492059 633326 492473
rect 136 491829 633326 492059
rect 0 491602 633326 491829
rect -2 491507 633326 491602
rect -2 491466 58 491507
rect -2 491427 122 491466
rect 136 491277 633326 491507
rect 0 489023 633326 491277
rect 136 488793 633326 489023
rect 0 488474 633326 488793
rect -2 488379 633326 488474
rect -2 488338 58 488379
rect -2 488299 122 488338
rect 136 488149 633326 488379
rect 0 487735 633326 488149
rect 136 487505 633326 487735
rect 0 487183 633326 487505
rect 136 486953 633326 487183
rect 0 485343 633326 486953
rect 136 485113 633326 485343
rect 0 484699 633326 485113
rect 136 484469 633326 484699
rect 0 484055 633326 484469
rect 136 483825 633326 484055
rect 0 483503 633326 483825
rect 136 483273 633326 483503
rect 0 478784 633326 483273
rect 136 478564 633326 478784
rect 0 476784 633326 478564
rect 136 476564 633326 476784
rect 0 432563 633326 476564
rect 0 417723 633571 432563
rect 0 370623 633326 417723
rect 136 370393 633326 370623
rect 0 368783 633326 370393
rect -2 368598 122 368633
rect -2 368553 58 368598
rect 136 368553 633326 368783
rect -2 368462 633326 368553
rect 0 368139 633326 368462
rect 136 367909 633326 368139
rect 0 366943 633326 367909
rect 136 366713 633326 366943
rect 0 366299 633326 366713
rect 136 366069 633326 366299
rect 0 365747 633326 366069
rect 136 365517 633326 365747
rect 0 365103 633326 365517
rect 136 364873 633326 365103
rect 0 364459 633326 364873
rect 136 364229 633326 364459
rect 0 363907 633326 364229
rect 136 363677 633326 363907
rect 0 361423 633326 363677
rect 136 361193 633326 361423
rect 0 360779 633326 361193
rect 136 360549 633326 360779
rect 0 360135 633326 360549
rect 136 359905 633326 360135
rect 0 359583 633326 359905
rect 136 359353 633326 359583
rect 0 357743 633326 359353
rect 136 357513 633326 357743
rect 0 357099 633326 357513
rect 136 356869 633326 357099
rect 0 356455 633326 356869
rect 136 356225 633326 356455
rect 0 355903 633326 356225
rect 136 355673 633326 355903
rect 0 349890 633326 355673
rect -2 349784 633326 349890
rect -2 349754 58 349784
rect -2 349704 122 349754
rect 136 349564 633326 349784
rect 0 348258 633326 349564
rect 0 348149 633328 348258
rect 0 347927 633190 348149
rect 633268 348122 633328 348149
rect 633206 348069 633328 348122
rect 0 347784 633326 347927
rect 136 347564 633326 347784
rect 0 346147 633326 347564
rect 0 345925 633190 346147
rect 0 344253 633326 345925
rect 0 344023 633190 344253
rect 0 343701 633326 344023
rect 0 343471 633190 343701
rect 0 343057 633326 343471
rect 0 342827 633190 343057
rect 0 342413 633326 342827
rect 0 342183 633190 342413
rect 0 340573 633326 342183
rect 0 340343 633190 340573
rect 0 340021 633326 340343
rect 0 339791 633190 340021
rect 0 339377 633326 339791
rect 0 339147 633190 339377
rect 0 338733 633326 339147
rect 0 338503 633190 338733
rect 633206 338542 633328 338583
rect 633268 338503 633328 338542
rect 0 338134 633328 338503
rect 0 336249 633326 338134
rect 0 336019 633190 336249
rect 0 335697 633326 336019
rect 0 335467 633190 335697
rect 0 335053 633326 335467
rect 0 334823 633190 335053
rect 633206 334870 633328 334903
rect 633268 334823 633328 334870
rect 0 334598 633328 334823
rect 0 334409 633326 334598
rect 0 334179 633190 334409
rect 0 333857 633326 334179
rect 0 333627 633190 333857
rect 0 333213 633326 333627
rect 0 332983 633190 333213
rect 0 332017 633326 332983
rect 0 331787 633190 332017
rect 0 331373 633326 331787
rect 0 331143 633190 331373
rect 0 329762 633326 331143
rect 0 329533 633328 329762
rect 0 329303 633190 329533
rect 633268 329490 633328 329533
rect 633206 329453 633328 329490
rect 0 327423 633326 329303
rect 136 327193 633326 327423
rect 0 325583 633326 327193
rect 136 325353 633326 325583
rect 0 324939 633326 325353
rect 136 324709 633326 324939
rect 0 323743 633326 324709
rect 136 323513 633326 323743
rect 0 323099 633326 323513
rect 136 322869 633326 323099
rect 0 322547 633326 322869
rect 136 322317 633326 322547
rect 0 322010 633326 322317
rect -2 321903 633326 322010
rect -2 321874 58 321903
rect -2 321823 122 321874
rect 136 321673 633326 321903
rect 0 321259 633326 321673
rect 136 321029 633326 321259
rect 0 320707 633326 321029
rect 136 320477 633326 320707
rect 0 318223 633326 320477
rect 136 317993 633326 318223
rect 0 317579 633326 317993
rect 136 317349 633326 317579
rect 0 316935 633326 317349
rect 136 316705 633326 316935
rect 0 316383 633326 316705
rect 136 316153 633326 316383
rect 0 314543 633326 316153
rect 136 314313 633326 314543
rect 0 313899 633326 314313
rect 136 313669 633326 313899
rect 0 313255 633326 313669
rect 136 313025 633326 313255
rect 0 312703 633326 313025
rect 136 312473 633326 312703
rect 0 306784 633326 312473
rect 136 306564 633326 306784
rect 0 304874 633326 306564
rect -2 304784 633326 304874
rect -2 304738 58 304784
rect -2 304704 122 304738
rect 136 304564 633326 304784
rect 0 303149 633326 304564
rect 0 302927 633190 303149
rect 0 301147 633326 302927
rect 0 300925 633190 301147
rect 0 299053 633326 300925
rect 0 298823 633190 299053
rect 0 298501 633326 298823
rect 0 298271 633190 298501
rect 0 297857 633326 298271
rect 0 297627 633190 297857
rect 0 297213 633326 297627
rect 0 296983 633190 297213
rect 0 295373 633326 296983
rect 0 295143 633190 295373
rect 0 294821 633326 295143
rect 0 294591 633190 294821
rect 0 294266 633326 294591
rect 0 294177 633328 294266
rect 0 293947 633190 294177
rect 633268 294130 633328 294177
rect 633206 294097 633328 294130
rect 0 293533 633326 293947
rect 0 293303 633190 293533
rect 0 291049 633326 293303
rect 0 290819 633190 291049
rect 0 290497 633326 290819
rect 0 290267 633190 290497
rect 0 289853 633326 290267
rect 0 289623 633190 289853
rect 0 289209 633326 289623
rect 0 288979 633190 289209
rect 0 288657 633326 288979
rect 0 288427 633190 288657
rect 0 288013 633326 288427
rect 0 287783 633190 288013
rect 633206 287814 633328 287863
rect 633268 287783 633328 287814
rect 0 287678 633328 287783
rect 0 286817 633326 287678
rect 0 286587 633190 286817
rect 0 286173 633326 286587
rect 0 285943 633190 286173
rect 0 284333 633326 285943
rect 0 284223 633190 284333
rect 136 284103 633190 284223
rect 136 283993 633326 284103
rect 0 282383 633326 283993
rect 136 282153 633326 282383
rect 0 281739 633326 282153
rect 136 281509 633326 281739
rect 0 280543 633326 281509
rect 136 280313 633326 280543
rect 0 279899 633326 280313
rect 136 279669 633326 279899
rect 0 279442 633326 279669
rect -2 279347 633326 279442
rect -2 279306 58 279347
rect -2 279267 122 279306
rect 136 279117 633326 279347
rect 0 278703 633326 279117
rect 136 278473 633326 278703
rect 0 278059 633326 278473
rect 136 277829 633326 278059
rect 0 277507 633326 277829
rect 136 277277 633326 277507
rect 0 275023 633326 277277
rect 136 274793 633326 275023
rect 0 274379 633326 274793
rect 136 274149 633326 274379
rect 0 273735 633326 274149
rect 136 273505 633326 273735
rect 0 273183 633326 273505
rect 136 272953 633326 273183
rect 0 271343 633326 272953
rect 136 271113 633326 271343
rect 0 270699 633326 271113
rect 136 270469 633326 270699
rect 0 270055 633326 270469
rect 136 269825 633326 270055
rect 0 269503 633326 269825
rect 136 269273 633326 269503
rect 0 263784 633326 269273
rect 136 263564 633326 263784
rect 0 261784 633326 263564
rect 136 261564 633326 261784
rect 0 258149 633326 261564
rect 0 257927 633190 258149
rect 0 256147 633326 257927
rect 0 255925 633190 256147
rect 0 254053 633326 255925
rect 0 253823 633190 254053
rect 0 253602 633326 253823
rect 0 253501 633328 253602
rect 0 253271 633190 253501
rect 633268 253466 633328 253501
rect 633206 253421 633328 253466
rect 0 252857 633326 253271
rect 0 252627 633190 252857
rect 0 252213 633326 252627
rect 0 251983 633190 252213
rect 0 250373 633326 251983
rect 0 250143 633190 250373
rect 0 249821 633326 250143
rect 0 249591 633190 249821
rect 0 249177 633326 249591
rect 0 248947 633190 249177
rect 0 248533 633326 248947
rect 0 248303 633190 248533
rect 0 246049 633326 248303
rect 0 245819 633190 246049
rect 0 245497 633326 245819
rect 0 245267 633190 245497
rect 0 244853 633326 245267
rect 0 244623 633190 244853
rect 0 244209 633326 244623
rect 0 243979 633190 244209
rect 633206 244022 633328 244059
rect 633268 243979 633328 244022
rect 0 243886 633328 243979
rect 0 243657 633326 243886
rect 0 243427 633190 243657
rect 0 243013 633326 243427
rect 0 242783 633190 243013
rect 0 241817 633326 242783
rect 0 241587 633190 241817
rect 0 241173 633326 241587
rect 0 241023 633190 241173
rect 136 240943 633190 241023
rect 136 240793 633326 240943
rect 0 239333 633326 240793
rect 0 239183 633190 239333
rect 136 239103 633190 239183
rect 136 238953 633326 239103
rect 0 238539 633326 238953
rect 136 238309 633326 238539
rect 0 237343 633326 238309
rect 136 237113 633326 237343
rect 0 236699 633326 237113
rect 136 236469 633326 236699
rect 0 236147 633326 236469
rect 136 235917 633326 236147
rect 0 235503 633326 235917
rect -2 235318 122 235353
rect -2 235273 58 235318
rect 136 235273 633326 235503
rect -2 235182 633326 235273
rect 0 234970 633326 235182
rect -2 234859 633326 234970
rect -2 234834 58 234859
rect -2 234779 122 234834
rect 136 234629 633326 234859
rect 0 234307 633326 234629
rect 136 234077 633326 234307
rect 0 231823 633326 234077
rect 136 231593 633326 231823
rect 0 231179 633326 231593
rect 136 230949 633326 231179
rect 0 230535 633326 230949
rect 136 230305 633326 230535
rect 0 230074 633326 230305
rect -2 229983 633326 230074
rect -2 229938 58 229983
rect -2 229903 122 229938
rect 136 229753 633326 229983
rect 0 228143 633326 229753
rect 136 227913 633326 228143
rect 0 227499 633326 227913
rect 136 227269 633326 227499
rect 0 226855 633326 227269
rect 136 226625 633326 226855
rect 0 226303 633326 226625
rect 136 226073 633326 226303
rect 0 220784 633326 226073
rect 136 220564 633326 220784
rect 0 218784 633326 220564
rect 136 218564 633326 218784
rect 0 213149 633326 218564
rect 0 212927 633190 213149
rect 0 211147 633326 212927
rect 0 210925 633190 211147
rect 633206 210974 633328 211005
rect 633268 210925 633328 210974
rect 0 210838 633328 210925
rect 0 209053 633326 210838
rect 0 208823 633190 209053
rect 0 208501 633326 208823
rect 0 208271 633190 208501
rect 0 207857 633326 208271
rect 0 207627 633190 207857
rect 0 207213 633326 207627
rect 0 206983 633190 207213
rect 0 205373 633326 206983
rect 0 205143 633190 205373
rect 0 204821 633326 205143
rect 0 204591 633190 204821
rect 0 204177 633326 204591
rect 0 203947 633190 204177
rect 0 203533 633326 203947
rect 0 203303 633190 203533
rect 0 201049 633326 203303
rect 0 200819 633190 201049
rect 0 200497 633326 200819
rect 0 200267 633190 200497
rect 0 199853 633326 200267
rect 0 199623 633190 199853
rect 0 199209 633326 199623
rect 0 198979 633190 199209
rect 633206 199006 633328 199059
rect 633268 198979 633328 199006
rect 0 198734 633328 198979
rect 0 198657 633326 198734
rect 0 198427 633190 198657
rect 0 198013 633326 198427
rect 0 197824 633190 198013
rect 136 197783 633190 197824
rect 136 197592 633326 197783
rect 0 196817 633326 197592
rect 0 196587 633190 196817
rect 0 196173 633326 196587
rect 0 195984 633190 196173
rect 136 195943 633190 195984
rect 136 195752 633326 195943
rect 0 195340 633326 195752
rect 136 195108 633326 195340
rect 0 194333 633326 195108
rect 0 194144 633190 194333
rect 136 194103 633190 194144
rect 136 193912 633326 194103
rect 0 193500 633326 193912
rect 136 193268 633326 193500
rect 0 192948 633326 193268
rect 136 192716 633326 192948
rect 0 192402 633326 192716
rect -2 192304 633326 192402
rect -2 192266 58 192304
rect -2 192224 122 192266
rect 136 192072 633326 192304
rect 0 191660 633326 192072
rect 136 191428 633326 191660
rect 0 191108 633326 191428
rect 136 190876 633326 191108
rect 0 188866 633326 190876
rect -2 188624 633326 188866
rect -2 188594 58 188624
rect -2 188544 122 188594
rect 136 188392 633326 188624
rect 0 187980 633326 188392
rect 136 187748 633326 187980
rect 0 187336 633326 187748
rect 136 187104 633326 187336
rect 0 186784 633326 187104
rect 136 186552 633326 186784
rect 0 184944 633326 186552
rect 136 184712 633326 184944
rect 0 184300 633326 184712
rect 136 184068 633326 184300
rect 0 183656 633326 184068
rect 136 183424 633326 183656
rect 0 183104 633326 183424
rect 136 182872 633326 183104
rect 0 177986 633326 182872
rect -2 177790 633326 177986
rect 0 177784 633326 177790
rect 136 177564 633326 177784
rect 0 175784 633326 177564
rect 136 175564 633326 175784
rect 0 168149 633326 175564
rect 0 167927 633190 168149
rect 0 166147 633326 167927
rect 0 165925 633190 166147
rect 0 163853 633326 165925
rect 0 163623 633190 163853
rect 0 163301 633326 163623
rect 0 163071 633190 163301
rect 0 162657 633326 163071
rect 0 162427 633190 162657
rect 0 162013 633326 162427
rect 0 161783 633190 162013
rect 0 160173 633326 161783
rect 0 159943 633190 160173
rect 0 159621 633326 159943
rect 0 159391 633190 159621
rect 633206 159430 633328 159471
rect 633268 159391 633328 159430
rect 0 159294 633328 159391
rect 0 158977 633326 159294
rect 0 158747 633190 158977
rect 0 158333 633326 158747
rect 0 158103 633190 158333
rect 0 155849 633326 158103
rect 0 155619 633190 155849
rect 0 155297 633326 155619
rect 0 155067 633190 155297
rect 0 154653 633326 155067
rect 0 154624 633190 154653
rect 136 154423 633190 154624
rect 136 154392 633326 154423
rect 0 154009 633326 154392
rect 0 153779 633190 154009
rect 0 153457 633326 153779
rect 0 153227 633190 153457
rect 0 152813 633326 153227
rect 0 152784 633190 152813
rect 136 152583 633190 152784
rect 136 152552 633326 152583
rect 0 152140 633326 152552
rect 136 151908 633326 152140
rect 0 151617 633326 151908
rect 0 151387 633190 151617
rect 0 150973 633326 151387
rect 0 150944 633190 150973
rect 136 150743 633190 150944
rect 136 150712 633326 150743
rect 0 150300 633326 150712
rect 136 150068 633326 150300
rect 0 149748 633326 150068
rect 136 149516 633326 149748
rect 0 149133 633326 149516
rect 0 149104 633190 149133
rect 136 148903 633190 149104
rect 136 148872 633326 148903
rect 0 148460 633326 148872
rect 136 148228 633326 148460
rect 0 147908 633326 148228
rect 136 147676 633326 147908
rect 0 145424 633326 147676
rect 136 145192 633326 145424
rect 0 144780 633326 145192
rect 136 144548 633326 144780
rect 0 144136 633326 144548
rect 136 143904 633326 144136
rect 0 143584 633326 143904
rect 136 143352 633326 143584
rect 0 141744 633326 143352
rect 136 141512 633326 141744
rect 0 141100 633326 141512
rect 136 140868 633326 141100
rect 0 140456 633326 140868
rect 136 140224 633326 140456
rect 0 139904 633326 140224
rect 136 139672 633326 139904
rect 0 135010 633326 139672
rect -2 134784 633326 135010
rect -2 134738 58 134784
rect -2 134704 122 134738
rect 136 134564 633326 134784
rect 0 132784 633326 134564
rect 136 132564 633326 132784
rect 0 123149 633326 132564
rect 0 122927 633190 123149
rect 0 121147 633326 122927
rect 0 120925 633190 121147
rect 0 118853 633326 120925
rect 0 118623 633190 118853
rect 0 118301 633326 118623
rect 0 118071 633190 118301
rect 0 117657 633326 118071
rect 0 117427 633190 117657
rect 0 117013 633326 117427
rect 0 116783 633190 117013
rect 0 115173 633326 116783
rect 0 114943 633190 115173
rect 0 114621 633326 114943
rect 0 114391 633190 114621
rect 0 113977 633326 114391
rect 0 113747 633190 113977
rect 0 113333 633326 113747
rect 0 113103 633190 113333
rect 0 110938 633326 113103
rect 0 110849 633328 110938
rect 0 110619 633190 110849
rect 633268 110802 633328 110849
rect 633206 110769 633328 110802
rect 0 110297 633326 110619
rect 0 110067 633190 110297
rect 0 109653 633326 110067
rect 0 109423 633190 109653
rect 0 109009 633326 109423
rect 0 108779 633190 109009
rect 0 108457 633326 108779
rect 0 108227 633190 108457
rect 0 107813 633326 108227
rect 0 107583 633190 107813
rect 0 106617 633326 107583
rect 0 106387 633190 106617
rect 0 105973 633326 106387
rect 0 105743 633190 105973
rect 0 104133 633326 105743
rect 0 103903 633190 104133
rect 0 78149 633326 103903
rect 0 77927 633190 78149
rect 0 76258 633326 77927
rect 0 76147 633328 76258
rect 0 75925 633190 76147
rect 633268 76122 633328 76147
rect 633206 76067 633328 76122
rect 0 73653 633326 75925
rect 0 73423 633190 73653
rect 0 73101 633326 73423
rect 0 72871 633190 73101
rect 0 72457 633326 72871
rect 0 72227 633190 72457
rect 633206 72254 633328 72307
rect 633268 72227 633328 72254
rect 0 72118 633328 72227
rect 0 71813 633326 72118
rect 0 71583 633190 71813
rect 0 69973 633326 71583
rect 0 69743 633190 69973
rect 0 69421 633326 69743
rect 0 69191 633190 69421
rect 0 68777 633326 69191
rect 0 68547 633190 68777
rect 633206 68582 633328 68627
rect 633268 68547 633328 68582
rect 0 68174 633328 68547
rect 0 68133 633326 68174
rect 0 67903 633190 68133
rect 0 65649 633326 67903
rect 0 65419 633190 65649
rect 0 65097 633326 65419
rect 0 64867 633190 65097
rect 0 64453 633326 64867
rect 0 64223 633190 64453
rect 0 63809 633326 64223
rect 0 63579 633190 63809
rect 0 63257 633326 63579
rect 0 63027 633190 63257
rect 0 62613 633326 63027
rect 0 62383 633190 62613
rect 0 61417 633326 62383
rect 0 61187 633190 61417
rect 0 60773 633326 61187
rect 0 60543 633190 60773
rect 0 58933 633326 60543
rect 0 58703 633190 58933
rect 0 53745 633326 58703
rect 136 53067 633326 53745
rect 0 8127 633326 53067
<< metal4 >>
rect 324 480 4324 952608
rect 4804 4960 8804 948128
rect 11050 480 12330 952608
rect 12970 480 14250 952608
rect 19050 480 20330 952608
rect 20970 480 22250 952608
rect 27050 480 28330 952608
rect 28970 480 30250 952608
rect 35050 480 36330 952608
rect 36970 480 38250 952608
rect 43050 480 44330 952608
rect 44970 480 46250 952608
rect 51050 480 52330 952608
rect 52970 480 54250 952608
rect 59050 480 60330 952608
rect 60970 480 62250 952608
rect 67050 480 68330 952608
rect 68970 480 70250 952608
rect 75050 480 76330 952608
rect 76970 480 78250 952608
rect 83050 480 84330 952608
rect 84970 480 86250 952608
rect 91050 709904 92330 952608
rect 92970 709904 94250 952608
rect 99050 709904 100330 952608
rect 100970 709904 102250 952608
rect 107050 709904 108330 952608
rect 108970 709904 110250 952608
rect 115050 709904 116330 952608
rect 116970 709904 118250 952608
rect 123050 709904 124330 952608
rect 124970 709904 126250 952608
rect 131050 709904 132330 952608
rect 132970 709904 134250 952608
rect 139050 709904 140330 952608
rect 140970 709904 142250 952608
rect 147050 709904 148330 952608
rect 148970 709904 150250 952608
rect 155050 709904 156330 952608
rect 156970 709904 158250 952608
rect 163050 709904 164330 952608
rect 164970 709904 166250 952608
rect 171050 709904 172330 952608
rect 172970 709904 174250 952608
rect 179050 709904 180330 952608
rect 180970 709904 182250 952608
rect 187050 709904 188330 952608
rect 188970 709904 190250 952608
rect 195050 709904 196330 952608
rect 196970 709904 198250 952608
rect 203050 709904 204330 952608
rect 204970 709904 206250 952608
rect 211050 709904 212330 952608
rect 212970 709904 214250 952608
rect 219050 709904 220330 952608
rect 220970 709904 222250 952608
rect 227050 709904 228330 952608
rect 228970 709904 230250 952608
rect 235050 709904 236330 952608
rect 236970 709904 238250 952608
rect 243050 709904 244330 952608
rect 244970 709904 246250 952608
rect 251050 709904 252330 952608
rect 252970 709904 254250 952608
rect 259050 709904 260330 952608
rect 260970 709904 262250 952608
rect 267050 709904 268330 952608
rect 268970 709904 270250 952608
rect 275050 709904 276330 952608
rect 276970 709904 278250 952608
rect 283050 709904 284330 952608
rect 284970 709904 286250 952608
rect 291050 709904 292330 952608
rect 292970 709904 294250 952608
rect 299050 709904 300330 952608
rect 300970 709904 302250 952608
rect 307050 709904 308330 952608
rect 308970 709904 310250 952608
rect 315050 709904 316330 952608
rect 316970 709904 318250 952608
rect 323050 709904 324330 952608
rect 324970 709904 326250 952608
rect 331050 709904 332330 952608
rect 332970 709904 334250 952608
rect 339050 709904 340330 952608
rect 340970 709904 342250 952608
rect 347050 709904 348330 952608
rect 348970 709904 350250 952608
rect 355050 709904 356330 952608
rect 356970 709904 358250 952608
rect 363050 709904 364330 952608
rect 364970 709904 366250 952608
rect 371050 709904 372330 952608
rect 372970 709904 374250 952608
rect 379050 709904 380330 952608
rect 380970 709904 382250 952608
rect 387050 709904 388330 952608
rect 388970 709904 390250 952608
rect 395050 709904 396330 952608
rect 396970 709904 398250 952608
rect 403050 709904 404330 952608
rect 404970 709904 406250 952608
rect 411050 709904 412330 952608
rect 412970 709904 414250 952608
rect 419050 709904 420330 952608
rect 420970 709904 422250 952608
rect 427050 709904 428330 952608
rect 428970 709904 430250 952608
rect 435050 709904 436330 952608
rect 436970 709904 438250 952608
rect 443050 709904 444330 952608
rect 444970 709904 446250 952608
rect 451050 709904 452330 952608
rect 452970 709904 454250 952608
rect 459050 709904 460330 952608
rect 460970 709904 462250 952608
rect 467050 709904 468330 952608
rect 468970 709904 470250 952608
rect 475050 709904 476330 952608
rect 476970 709904 478250 952608
rect 483050 709904 484330 952608
rect 484970 709904 486250 952608
rect 491050 709904 492330 952608
rect 492970 709904 494250 952608
rect 499050 709904 500330 952608
rect 500970 709904 502250 952608
rect 507050 709904 508330 952608
rect 508970 709904 510250 952608
rect 515050 709904 516330 952608
rect 516970 709904 518250 952608
rect 523050 709904 524330 952608
rect 524970 709904 526250 952608
rect 531050 709904 532330 952608
rect 532970 709904 534250 952608
rect 539050 709904 540330 952608
rect 540970 709904 542250 952608
rect 547050 709904 548330 952608
rect 548970 709904 550250 952608
rect 555050 709904 556330 952608
rect 556970 709904 558250 952608
rect 563050 709904 564330 952608
rect 564970 709904 566250 952608
rect 571050 709904 572330 952608
rect 572970 709904 574250 952608
rect 579050 709904 580330 952608
rect 580970 709904 582250 952608
rect 587050 709904 588330 952608
rect 588970 709904 590250 952608
rect 595050 709904 596330 952608
rect 596970 709904 598250 952608
rect 603050 709904 604330 952608
rect 604970 709904 606250 952608
rect 91050 480 92330 389968
rect 92970 480 94250 389968
rect 99050 480 100330 389968
rect 100970 480 102250 389968
rect 107050 480 108330 389968
rect 108970 480 110250 389968
rect 115050 480 116330 389968
rect 116970 480 118250 389968
rect 123050 480 124330 389968
rect 124970 480 126250 389968
rect 131050 480 132330 389968
rect 132970 480 134250 389968
rect 139050 480 140330 389968
rect 140970 480 142250 389968
rect 147050 480 148330 389968
rect 148970 480 150250 389968
rect 155050 480 156330 389968
rect 156970 480 158250 389968
rect 163050 480 164330 389968
rect 164970 480 166250 389968
rect 171050 480 172330 389968
rect 172970 480 174250 389968
rect 179050 480 180330 389968
rect 180970 480 182250 389968
rect 187050 480 188330 389968
rect 188970 480 190250 389968
rect 195050 480 196330 389968
rect 196970 480 198250 389968
rect 203050 480 204330 389968
rect 204970 480 206250 389968
rect 211050 480 212330 389968
rect 212970 480 214250 389968
rect 219050 480 220330 389968
rect 220970 480 222250 389968
rect 227050 480 228330 389968
rect 228970 480 230250 389968
rect 235050 480 236330 389968
rect 236970 480 238250 389968
rect 243050 480 244330 389968
rect 244970 480 246250 389968
rect 251050 480 252330 389968
rect 252970 480 254250 389968
rect 259050 480 260330 389968
rect 260970 480 262250 389968
rect 267050 480 268330 389968
rect 268970 480 270250 389968
rect 275050 480 276330 389968
rect 276970 480 278250 389968
rect 283050 480 284330 389968
rect 284970 480 286250 389968
rect 291050 480 292330 389968
rect 292970 480 294250 389968
rect 299050 480 300330 389968
rect 300970 480 302250 389968
rect 307050 480 308330 389968
rect 308970 480 310250 389968
rect 315050 480 316330 389968
rect 316970 480 318250 389968
rect 323050 480 324330 389968
rect 324970 480 326250 389968
rect 331050 480 332330 389968
rect 332970 480 334250 389968
rect 339050 480 340330 389968
rect 340970 480 342250 389968
rect 347050 480 348330 389968
rect 348970 480 350250 389968
rect 355050 480 356330 389968
rect 356970 480 358250 389968
rect 363050 480 364330 389968
rect 364970 480 366250 389968
rect 371050 480 372330 389968
rect 372970 480 374250 389968
rect 379050 480 380330 389968
rect 380970 480 382250 389968
rect 387050 480 388330 389968
rect 388970 480 390250 389968
rect 395050 480 396330 389968
rect 396970 480 398250 389968
rect 403050 480 404330 389968
rect 404970 480 406250 389968
rect 411050 480 412330 389968
rect 412970 480 414250 389968
rect 419050 480 420330 389968
rect 420970 480 422250 389968
rect 427050 480 428330 389968
rect 428970 480 430250 389968
rect 435050 480 436330 389968
rect 436970 480 438250 389968
rect 443050 480 444330 389968
rect 444970 480 446250 389968
rect 451050 480 452330 389968
rect 452970 480 454250 389968
rect 459050 480 460330 389968
rect 460970 480 462250 389968
rect 467050 480 468330 389968
rect 468970 480 470250 389968
rect 475050 480 476330 389968
rect 476970 480 478250 389968
rect 483050 480 484330 389968
rect 484970 480 486250 389968
rect 491050 480 492330 389968
rect 492970 480 494250 389968
rect 499050 480 500330 389968
rect 500970 480 502250 389968
rect 507050 480 508330 389968
rect 508970 480 510250 389968
rect 515050 480 516330 389968
rect 516970 480 518250 389968
rect 523050 480 524330 389968
rect 524970 480 526250 389968
rect 531050 480 532330 389968
rect 532970 480 534250 389968
rect 539050 480 540330 389968
rect 540970 480 542250 389968
rect 547050 480 548330 389968
rect 548970 480 550250 389968
rect 555050 480 556330 389968
rect 556970 480 558250 389968
rect 563050 480 564330 389968
rect 564970 480 566250 389968
rect 571050 480 572330 389968
rect 572970 480 574250 389968
rect 579050 480 580330 389968
rect 580970 480 582250 389968
rect 587050 480 588330 389968
rect 588970 480 590250 389968
rect 595050 480 596330 389968
rect 596970 480 598250 389968
rect 603050 480 604330 389968
rect 604970 480 606250 389968
rect 611050 480 612330 952608
rect 612970 480 614250 952608
rect 619050 480 620330 952608
rect 620970 480 622250 952608
rect 624524 4960 628524 948128
rect 629004 480 633004 952608
<< obsm4 >>
rect 91794 390048 610970 707744
rect 92410 63411 92890 390048
rect 94330 63411 98970 390048
rect 100410 63411 100890 390048
rect 102330 63411 106970 390048
rect 108410 63411 108890 390048
rect 110330 63411 114970 390048
rect 116410 63411 116890 390048
rect 118330 63411 122970 390048
rect 124410 63411 124890 390048
rect 126330 63411 130970 390048
rect 132410 63411 132890 390048
rect 134330 63411 138970 390048
rect 140410 63411 140890 390048
rect 142330 63411 146970 390048
rect 148410 63411 148890 390048
rect 150330 63411 154970 390048
rect 156410 63411 156890 390048
rect 158330 63411 162970 390048
rect 164410 63411 164890 390048
rect 166330 63411 170970 390048
rect 172410 63411 172890 390048
rect 174330 63411 178970 390048
rect 180410 63411 180890 390048
rect 182330 63411 186970 390048
rect 188410 63411 188890 390048
rect 190330 63411 194970 390048
rect 196410 63411 196890 390048
rect 198330 63411 202970 390048
rect 204410 63411 204890 390048
rect 206330 63411 210970 390048
rect 212410 63411 212890 390048
rect 214330 63411 218970 390048
rect 220410 63411 220890 390048
rect 222330 63411 226970 390048
rect 228410 63411 228890 390048
rect 230330 63411 234970 390048
rect 236410 63411 236890 390048
rect 238330 63411 242970 390048
rect 244410 63411 244890 390048
rect 246330 63411 250970 390048
rect 252410 63411 252890 390048
rect 254330 63411 258970 390048
rect 260410 63411 260890 390048
rect 262330 63411 266970 390048
rect 268410 63411 268890 390048
rect 270330 63411 274970 390048
rect 276410 63411 276890 390048
rect 278330 63411 282970 390048
rect 284410 63411 284890 390048
rect 286330 63411 290970 390048
rect 292410 63411 292890 390048
rect 294330 63411 298970 390048
rect 300410 63411 300890 390048
rect 302330 63411 306970 390048
rect 308410 63411 308890 390048
rect 310330 63411 314970 390048
rect 316410 63411 316890 390048
rect 318330 63411 322970 390048
rect 324410 63411 324890 390048
rect 326330 63411 330970 390048
rect 332410 63411 332890 390048
rect 334330 63411 338970 390048
rect 340410 63411 340890 390048
rect 342330 63411 346970 390048
rect 348410 63411 348890 390048
rect 350330 63411 354970 390048
rect 356410 63411 356890 390048
rect 358330 63411 362970 390048
rect 364410 63411 364890 390048
rect 366330 63411 370970 390048
rect 372410 63411 372890 390048
rect 374330 63411 378970 390048
rect 380410 63411 380890 390048
rect 382330 63411 386970 390048
rect 388410 63411 388890 390048
rect 390330 63411 394970 390048
rect 396410 63411 396890 390048
rect 398330 63411 402970 390048
rect 404410 63411 404890 390048
rect 406330 63411 410970 390048
rect 412410 63411 412890 390048
rect 414330 63411 418970 390048
rect 420410 63411 420890 390048
rect 422330 63411 426970 390048
rect 428410 63411 428890 390048
rect 430330 63411 434970 390048
rect 436410 63411 436890 390048
rect 438330 63411 442970 390048
rect 444410 63411 444890 390048
rect 446330 63411 450970 390048
rect 452410 63411 452890 390048
rect 454330 63411 458970 390048
rect 460410 63411 460890 390048
rect 462330 63411 466970 390048
rect 468410 63411 468890 390048
rect 470330 63411 474970 390048
rect 476410 63411 476890 390048
rect 478330 63411 482970 390048
rect 484410 63411 484890 390048
rect 486330 63411 490970 390048
rect 492410 63411 492890 390048
rect 494330 63411 498970 390048
rect 500410 63411 500890 390048
rect 502330 63411 506970 390048
rect 508410 63411 508890 390048
rect 510330 63411 514970 390048
rect 516410 63411 516890 390048
rect 518330 63411 522970 390048
rect 524410 63411 524890 390048
rect 526330 63411 530970 390048
rect 532410 63411 532890 390048
rect 534330 63411 538970 390048
rect 540410 63411 540890 390048
rect 542330 63411 546970 390048
rect 548410 63411 548890 390048
rect 550330 63411 554970 390048
rect 556410 63411 556890 390048
rect 558330 63411 562970 390048
rect 564410 63411 564890 390048
rect 566330 63411 570970 390048
rect 572410 63411 572890 390048
rect 574330 63411 578970 390048
rect 580410 63411 580890 390048
rect 582330 63411 586970 390048
rect 588410 63411 588890 390048
rect 590330 63411 594970 390048
rect 596410 63411 596890 390048
rect 598330 63411 602970 390048
rect 604410 63411 604890 390048
rect 606330 63411 610970 390048
rect 612410 63411 612890 707744
rect 614330 63411 618970 707744
rect 620410 63411 620890 707744
rect 622330 63411 624437 707744
<< metal5 >>
rect 324 948608 633004 952608
rect 4804 944128 628524 948128
rect 324 942006 633004 943286
rect 324 940086 633004 941366
rect 324 934006 633004 935286
rect 324 932086 633004 933366
rect 324 926006 633004 927286
rect 324 924086 633004 925366
rect 324 918006 633004 919286
rect 324 916086 633004 917366
rect 324 910006 633004 911286
rect 324 908086 633004 909366
rect 324 902006 633004 903286
rect 324 900086 633004 901366
rect 324 894006 633004 895286
rect 324 892086 633004 893366
rect 324 886006 633004 887286
rect 324 884086 633004 885366
rect 324 878006 633004 879286
rect 324 876086 633004 877366
rect 324 870006 633004 871286
rect 324 868086 633004 869366
rect 324 862006 633004 863286
rect 324 860086 633004 861366
rect 324 854006 633004 855286
rect 324 852086 633004 853366
rect 324 846006 633004 847286
rect 324 844086 633004 845366
rect 324 838006 633004 839286
rect 324 836086 633004 837366
rect 324 830006 633004 831286
rect 324 828086 633004 829366
rect 324 822006 633004 823286
rect 324 820086 633004 821366
rect 324 814006 633004 815286
rect 324 812086 633004 813366
rect 324 806006 633004 807286
rect 324 804086 633004 805366
rect 324 798006 633004 799286
rect 324 796086 633004 797366
rect 324 790006 633004 791286
rect 324 788086 633004 789366
rect 324 782006 633004 783286
rect 324 780086 633004 781366
rect 324 774006 633004 775286
rect 324 772086 633004 773366
rect 324 766006 633004 767286
rect 324 764086 633004 765366
rect 324 758006 633004 759286
rect 324 756086 633004 757366
rect 324 750006 633004 751286
rect 324 748086 633004 749366
rect 324 742006 633004 743286
rect 324 740086 633004 741366
rect 324 734006 633004 735286
rect 324 732086 633004 733366
rect 324 726006 633004 727286
rect 324 724086 633004 725366
rect 324 718006 633004 719286
rect 324 716086 633004 717366
rect 324 710006 633004 711286
rect 324 708086 633004 709366
rect 324 702006 633004 703286
rect 324 700086 633004 701366
rect 324 694006 633004 695286
rect 324 692086 633004 693366
rect 324 686006 633004 687286
rect 324 684086 633004 685366
rect 324 678006 633004 679286
rect 324 676086 633004 677366
rect 324 670006 633004 671286
rect 324 668086 633004 669366
rect 324 662006 633004 663286
rect 324 660086 633004 661366
rect 324 654006 633004 655286
rect 324 652086 633004 653366
rect 324 646006 633004 647286
rect 324 644086 633004 645366
rect 324 638006 633004 639286
rect 324 636086 633004 637366
rect 324 630006 633004 631286
rect 324 628086 633004 629366
rect 324 622006 633004 623286
rect 324 620086 633004 621366
rect 324 614006 633004 615286
rect 324 612086 633004 613366
rect 324 606006 633004 607286
rect 324 604086 633004 605366
rect 324 598006 633004 599286
rect 324 596086 633004 597366
rect 324 590006 633004 591286
rect 324 588086 633004 589366
rect 324 582006 633004 583286
rect 324 580086 633004 581366
rect 324 574006 633004 575286
rect 324 572086 633004 573366
rect 324 566006 633004 567286
rect 324 564086 633004 565366
rect 324 558006 633004 559286
rect 324 556086 633004 557366
rect 324 550006 633004 551286
rect 324 548086 633004 549366
rect 324 542006 139548 543286
rect 324 540086 139548 541366
rect 433660 542006 633004 543286
rect 433660 540086 633004 541366
rect 324 534006 139548 535286
rect 324 532086 139548 533366
rect 433660 534006 633004 535286
rect 433660 532086 633004 533366
rect 324 526006 139548 527286
rect 324 524086 139548 525366
rect 433660 526006 633004 527286
rect 433660 524086 633004 525366
rect 324 518006 139548 519286
rect 324 516086 139548 517366
rect 433660 518006 633004 519286
rect 433660 516086 633004 517366
rect 324 510006 139548 511286
rect 324 508086 139548 509366
rect 433660 510006 633004 511286
rect 433660 508086 633004 509366
rect 324 502006 139548 503286
rect 324 500086 139548 501366
rect 433660 502006 633004 503286
rect 433660 500086 633004 501366
rect 324 494006 139548 495286
rect 324 492086 139548 493366
rect 433660 494006 633004 495286
rect 433660 492086 633004 493366
rect 324 486006 139548 487286
rect 324 484086 139548 485366
rect 433660 486006 633004 487286
rect 433660 484086 633004 485366
rect 324 478006 139548 479286
rect 324 476086 139548 477366
rect 433660 478006 633004 479286
rect 433660 476086 633004 477366
rect 324 470006 139548 471286
rect 324 468086 139548 469366
rect 433660 470006 633004 471286
rect 433660 468086 633004 469366
rect 324 462006 139548 463286
rect 324 460086 139548 461366
rect 433660 462006 633004 463286
rect 433660 460086 633004 461366
rect 324 454006 139548 455286
rect 324 452086 139548 453366
rect 433660 454006 633004 455286
rect 433660 452086 633004 453366
rect 324 446006 633004 447286
rect 324 444086 633004 445366
rect 324 438006 633004 439286
rect 324 436086 633004 437366
rect 324 430006 633004 431286
rect 324 428086 633004 429366
rect 324 422006 633004 423286
rect 324 420086 633004 421366
rect 324 414006 633004 415286
rect 324 412086 633004 413366
rect 324 406006 633004 407286
rect 324 404086 633004 405366
rect 324 398006 633004 399286
rect 324 396086 633004 397366
rect 324 390006 633004 391286
rect 324 388086 633004 389366
rect 324 382006 633004 383286
rect 324 380086 633004 381366
rect 324 374006 633004 375286
rect 324 372086 633004 373366
rect 324 366006 633004 367286
rect 324 364086 633004 365366
rect 324 358006 633004 359286
rect 324 356086 633004 357366
rect 324 350006 633004 351286
rect 324 348086 633004 349366
rect 324 342006 633004 343286
rect 324 340086 633004 341366
rect 324 334006 633004 335286
rect 324 332086 633004 333366
rect 324 326006 633004 327286
rect 324 324086 633004 325366
rect 324 318006 633004 319286
rect 324 316086 633004 317366
rect 324 310006 633004 311286
rect 324 308086 633004 309366
rect 324 302006 633004 303286
rect 324 300086 633004 301366
rect 324 294006 633004 295286
rect 324 292086 633004 293366
rect 324 286006 633004 287286
rect 324 284086 633004 285366
rect 324 278006 633004 279286
rect 324 276086 633004 277366
rect 324 270006 633004 271286
rect 324 268086 633004 269366
rect 324 262006 633004 263286
rect 324 260086 633004 261366
rect 324 254006 633004 255286
rect 324 252086 633004 253366
rect 324 246006 633004 247286
rect 324 244086 633004 245366
rect 324 238006 633004 239286
rect 324 236086 633004 237366
rect 324 230006 633004 231286
rect 324 228086 633004 229366
rect 324 222006 633004 223286
rect 324 220086 633004 221366
rect 324 214006 633004 215286
rect 324 212086 633004 213366
rect 324 206006 633004 207286
rect 324 204086 633004 205366
rect 324 198006 633004 199286
rect 324 196086 633004 197366
rect 324 190006 633004 191286
rect 324 188086 633004 189366
rect 324 182006 633004 183286
rect 324 180086 633004 181366
rect 324 174006 633004 175286
rect 324 172086 633004 173366
rect 324 166006 633004 167286
rect 324 164086 633004 165366
rect 324 158006 633004 159286
rect 324 156086 633004 157366
rect 324 150006 633004 151286
rect 324 148086 633004 149366
rect 324 142006 633004 143286
rect 324 140086 633004 141366
rect 324 134006 633004 135286
rect 324 132086 633004 133366
rect 324 126006 633004 127286
rect 324 124086 633004 125366
rect 324 118006 633004 119286
rect 324 116086 633004 117366
rect 324 110006 633004 111286
rect 324 108086 633004 109366
rect 324 102006 633004 103286
rect 324 100086 633004 101366
rect 324 94006 633004 95286
rect 324 92086 633004 93366
rect 324 86006 633004 87286
rect 324 84086 633004 85366
rect 324 78006 633004 79286
rect 324 76086 633004 77366
rect 324 70006 633004 71286
rect 324 68086 633004 69366
rect 324 62006 633004 63286
rect 324 60086 633004 61366
rect 324 54006 633004 55286
rect 324 52086 633004 53366
rect 324 46006 633004 47286
rect 324 44086 633004 45366
rect 324 38006 633004 39286
rect 324 36086 633004 37366
rect 324 30006 633004 31286
rect 324 28086 633004 29366
rect 324 22006 633004 23286
rect 324 20086 633004 21366
rect 324 14006 633004 15286
rect 324 12086 633004 13366
rect 4804 4960 628524 8960
rect 324 480 633004 4480
<< obsm5 >>
rect 91056 703606 608928 706506
rect 91056 695606 608928 699766
rect 91056 687606 608928 691766
rect 91056 679606 608928 683766
rect 91056 671606 608928 675766
rect 91056 663606 608928 667766
rect 91056 655606 608928 659766
rect 91056 647606 608928 651766
rect 91056 639606 608928 643766
rect 91056 631606 608928 635766
rect 91056 623606 608928 627766
rect 91056 615606 608928 619766
rect 91056 607606 608928 611766
rect 91056 599606 608928 603766
rect 91056 591606 608928 595766
rect 91056 583606 608928 587766
rect 91056 575606 608928 579766
rect 91056 567606 608928 571766
rect 91056 559606 608928 563766
rect 91056 551606 608928 555766
rect 91056 543606 608928 547766
rect 139868 539766 433340 543606
rect 91056 535606 608928 539766
rect 139868 531766 433340 535606
rect 91056 527606 608928 531766
rect 139868 523766 433340 527606
rect 91056 519606 608928 523766
rect 139868 515766 433340 519606
rect 91056 511606 608928 515766
rect 139868 507766 433340 511606
rect 91056 503606 608928 507766
rect 139868 499766 433340 503606
rect 91056 495606 608928 499766
rect 139868 491766 433340 495606
rect 91056 487606 608928 491766
rect 139868 483766 433340 487606
rect 91056 479606 608928 483766
rect 139868 475766 433340 479606
rect 91056 471606 608928 475766
rect 139868 467766 433340 471606
rect 91056 463606 608928 467766
rect 139868 459766 433340 463606
rect 91056 455606 608928 459766
rect 139868 451766 433340 455606
rect 91056 447606 608928 451766
rect 91056 439606 608928 443766
rect 91056 431606 608928 435766
rect 91056 423606 608928 427766
rect 91056 415606 608928 419766
rect 91056 407606 608928 411766
rect 91056 399606 608928 403766
rect 91056 392866 608928 395766
<< labels >>
rlabel metal3 s 633270 61267 633750 61337 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 633270 644467 633750 644537 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 633270 689467 633750 689537 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 633270 734467 633750 734537 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 633270 823667 633750 823737 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 633270 912867 633750 912937 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 596396 953270 596452 953750 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 494596 953270 494652 953750 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 443196 953270 443252 953750 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 354196 953270 354252 953750 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 252396 953270 252452 953750 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 633270 106467 633750 106537 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 200796 953270 200852 953750 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 149396 953270 149452 953750 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 97996 953270 98052 953750 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 46596 953270 46652 953750 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -424 924589 56 924659 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -424 754789 56 754859 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -424 711589 56 711659 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -424 668389 56 668459 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -424 625189 56 625259 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s -424 581989 56 582059 4 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 633270 151467 633750 151537 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s -424 538789 56 538859 4 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s -424 495589 56 495659 4 analog_io[31]
port 25 nsew signal bidirectional
rlabel metal3 s -424 367989 56 368059 4 analog_io[32]
port 26 nsew signal bidirectional
rlabel metal3 s -424 324789 56 324859 4 analog_io[33]
port 27 nsew signal bidirectional
rlabel metal3 s -424 281589 56 281659 4 analog_io[34]
port 28 nsew signal bidirectional
rlabel metal3 s -424 238389 56 238459 4 analog_io[35]
port 29 nsew signal bidirectional
rlabel metal3 s -424 195188 56 195260 4 analog_io[36]
port 30 nsew signal bidirectional
rlabel metal3 s -424 151988 56 152060 4 analog_io[37]
port 31 nsew signal bidirectional
rlabel metal2 s 147674 -424 147730 56 8 analog_io[38]
port 32 nsew signal bidirectional
rlabel metal2 s 256274 -424 256330 56 8 analog_io[39]
port 33 nsew signal bidirectional
rlabel metal3 s 633270 196667 633750 196737 6 analog_io[3]
port 34 nsew signal bidirectional
rlabel metal2 s 311074 -424 311130 56 8 analog_io[40]
port 35 nsew signal bidirectional
rlabel metal2 s 365874 -424 365930 56 8 analog_io[41]
port 36 nsew signal bidirectional
rlabel metal2 s 420674 -424 420730 56 8 analog_io[42]
port 37 nsew signal bidirectional
rlabel metal2 s 475474 -424 475530 56 8 analog_io[43]
port 38 nsew signal bidirectional
rlabel metal3 s 633270 241667 633750 241737 6 analog_io[4]
port 39 nsew signal bidirectional
rlabel metal3 s 633270 286667 633750 286737 6 analog_io[5]
port 40 nsew signal bidirectional
rlabel metal3 s 633270 331867 633750 331937 6 analog_io[6]
port 41 nsew signal bidirectional
rlabel metal3 s 633270 509067 633750 509137 6 analog_io[7]
port 42 nsew signal bidirectional
rlabel metal3 s 633270 554267 633750 554337 6 analog_io[8]
port 43 nsew signal bidirectional
rlabel metal3 s 633270 599267 633750 599337 6 analog_io[9]
port 44 nsew signal bidirectional
rlabel metal3 s 633270 63107 633750 63177 6 analog_noesd_io[0]
port 45 nsew signal bidirectional
rlabel metal3 s 633270 646307 633750 646377 6 analog_noesd_io[10]
port 46 nsew signal bidirectional
rlabel metal3 s 633270 691307 633750 691377 6 analog_noesd_io[11]
port 47 nsew signal bidirectional
rlabel metal3 s 633270 736307 633750 736377 6 analog_noesd_io[12]
port 48 nsew signal bidirectional
rlabel metal3 s 633270 825507 633750 825577 6 analog_noesd_io[13]
port 49 nsew signal bidirectional
rlabel metal3 s 633270 914707 633750 914777 6 analog_noesd_io[14]
port 50 nsew signal bidirectional
rlabel metal2 s 594556 953270 594612 953750 6 analog_noesd_io[15]
port 51 nsew signal bidirectional
rlabel metal2 s 492756 953270 492812 953750 6 analog_noesd_io[16]
port 52 nsew signal bidirectional
rlabel metal2 s 441356 953270 441412 953750 6 analog_noesd_io[17]
port 53 nsew signal bidirectional
rlabel metal2 s 352356 953270 352412 953750 6 analog_noesd_io[18]
port 54 nsew signal bidirectional
rlabel metal2 s 250556 953270 250612 953750 6 analog_noesd_io[19]
port 55 nsew signal bidirectional
rlabel metal3 s 633270 108307 633750 108377 6 analog_noesd_io[1]
port 56 nsew signal bidirectional
rlabel metal2 s 198956 953270 199012 953750 6 analog_noesd_io[20]
port 57 nsew signal bidirectional
rlabel metal2 s 147556 953270 147612 953750 6 analog_noesd_io[21]
port 58 nsew signal bidirectional
rlabel metal2 s 96156 953270 96212 953750 6 analog_noesd_io[22]
port 59 nsew signal bidirectional
rlabel metal2 s 44756 953270 44812 953750 6 analog_noesd_io[23]
port 60 nsew signal bidirectional
rlabel metal3 s -424 922749 56 922819 4 analog_noesd_io[24]
port 61 nsew signal bidirectional
rlabel metal3 s -424 752949 56 753019 4 analog_noesd_io[25]
port 62 nsew signal bidirectional
rlabel metal3 s -424 709749 56 709819 4 analog_noesd_io[26]
port 63 nsew signal bidirectional
rlabel metal3 s -424 666549 56 666619 4 analog_noesd_io[27]
port 64 nsew signal bidirectional
rlabel metal3 s -424 623349 56 623419 4 analog_noesd_io[28]
port 65 nsew signal bidirectional
rlabel metal3 s -424 580149 56 580219 4 analog_noesd_io[29]
port 66 nsew signal bidirectional
rlabel metal3 s 633270 153307 633750 153377 6 analog_noesd_io[2]
port 67 nsew signal bidirectional
rlabel metal3 s -424 536949 56 537019 4 analog_noesd_io[30]
port 68 nsew signal bidirectional
rlabel metal3 s -424 493749 56 493819 4 analog_noesd_io[31]
port 69 nsew signal bidirectional
rlabel metal3 s -424 366149 56 366219 4 analog_noesd_io[32]
port 70 nsew signal bidirectional
rlabel metal3 s -424 322949 56 323019 4 analog_noesd_io[33]
port 71 nsew signal bidirectional
rlabel metal3 s -424 279749 56 279819 4 analog_noesd_io[34]
port 72 nsew signal bidirectional
rlabel metal3 s -424 236549 56 236619 4 analog_noesd_io[35]
port 73 nsew signal bidirectional
rlabel metal3 s -424 193348 56 193420 4 analog_noesd_io[36]
port 74 nsew signal bidirectional
rlabel metal3 s -424 150148 56 150220 4 analog_noesd_io[37]
port 75 nsew signal bidirectional
rlabel metal2 s 149514 -424 149570 56 8 analog_noesd_io[38]
port 76 nsew signal bidirectional
rlabel metal2 s 258114 -424 258170 56 8 analog_noesd_io[39]
port 77 nsew signal bidirectional
rlabel metal3 s 633270 198507 633750 198577 6 analog_noesd_io[3]
port 78 nsew signal bidirectional
rlabel metal2 s 312914 -424 312970 56 8 analog_noesd_io[40]
port 79 nsew signal bidirectional
rlabel metal2 s 367714 -424 367770 56 8 analog_noesd_io[41]
port 80 nsew signal bidirectional
rlabel metal2 s 422514 -424 422570 56 8 analog_noesd_io[42]
port 81 nsew signal bidirectional
rlabel metal2 s 477314 -424 477370 56 8 analog_noesd_io[43]
port 82 nsew signal bidirectional
rlabel metal3 s 633270 243507 633750 243577 6 analog_noesd_io[4]
port 83 nsew signal bidirectional
rlabel metal3 s 633270 288507 633750 288577 6 analog_noesd_io[5]
port 84 nsew signal bidirectional
rlabel metal3 s 633270 333707 633750 333777 6 analog_noesd_io[6]
port 85 nsew signal bidirectional
rlabel metal3 s 633270 510907 633750 510977 6 analog_noesd_io[7]
port 86 nsew signal bidirectional
rlabel metal3 s 633270 556107 633750 556177 6 analog_noesd_io[8]
port 87 nsew signal bidirectional
rlabel metal3 s 633270 601107 633750 601177 6 analog_noesd_io[9]
port 88 nsew signal bidirectional
rlabel metal3 s 633270 63659 633750 63729 6 gpio_analog_en[0]
port 89 nsew signal output
rlabel metal3 s 633270 646859 633750 646929 6 gpio_analog_en[10]
port 90 nsew signal output
rlabel metal3 s 633270 691859 633750 691929 6 gpio_analog_en[11]
port 91 nsew signal output
rlabel metal3 s 633270 736859 633750 736929 6 gpio_analog_en[12]
port 92 nsew signal output
rlabel metal3 s 633270 826059 633750 826129 6 gpio_analog_en[13]
port 93 nsew signal output
rlabel metal3 s 633270 915259 633750 915329 6 gpio_analog_en[14]
port 94 nsew signal output
rlabel metal2 s 594004 953270 594060 953750 6 gpio_analog_en[15]
port 95 nsew signal output
rlabel metal2 s 492204 953270 492260 953750 6 gpio_analog_en[16]
port 96 nsew signal output
rlabel metal2 s 440804 953270 440860 953750 6 gpio_analog_en[17]
port 97 nsew signal output
rlabel metal2 s 351804 953270 351860 953750 6 gpio_analog_en[18]
port 98 nsew signal output
rlabel metal2 s 250004 953270 250060 953750 6 gpio_analog_en[19]
port 99 nsew signal output
rlabel metal3 s 633270 108859 633750 108929 6 gpio_analog_en[1]
port 100 nsew signal output
rlabel metal2 s 198404 953270 198460 953750 6 gpio_analog_en[20]
port 101 nsew signal output
rlabel metal2 s 147004 953270 147060 953750 6 gpio_analog_en[21]
port 102 nsew signal output
rlabel metal2 s 95604 953270 95660 953750 6 gpio_analog_en[22]
port 103 nsew signal output
rlabel metal2 s 44204 953270 44260 953750 6 gpio_analog_en[23]
port 104 nsew signal output
rlabel metal3 s -424 922197 56 922267 4 gpio_analog_en[24]
port 105 nsew signal output
rlabel metal3 s -424 752397 56 752467 4 gpio_analog_en[25]
port 106 nsew signal output
rlabel metal3 s -424 709197 56 709267 4 gpio_analog_en[26]
port 107 nsew signal output
rlabel metal3 s -424 665997 56 666067 4 gpio_analog_en[27]
port 108 nsew signal output
rlabel metal3 s -424 622797 56 622867 4 gpio_analog_en[28]
port 109 nsew signal output
rlabel metal3 s -424 579597 56 579667 4 gpio_analog_en[29]
port 110 nsew signal output
rlabel metal3 s 633270 153859 633750 153929 6 gpio_analog_en[2]
port 111 nsew signal output
rlabel metal3 s -424 536397 56 536467 4 gpio_analog_en[30]
port 112 nsew signal output
rlabel metal3 s -424 493197 56 493267 4 gpio_analog_en[31]
port 113 nsew signal output
rlabel metal3 s -424 365597 56 365667 4 gpio_analog_en[32]
port 114 nsew signal output
rlabel metal3 s -424 322397 56 322467 4 gpio_analog_en[33]
port 115 nsew signal output
rlabel metal3 s -424 279197 56 279267 4 gpio_analog_en[34]
port 116 nsew signal output
rlabel metal3 s -424 235997 56 236067 4 gpio_analog_en[35]
port 117 nsew signal output
rlabel metal3 s -424 192796 56 192868 4 gpio_analog_en[36]
port 118 nsew signal output
rlabel metal3 s -424 149596 56 149668 4 gpio_analog_en[37]
port 119 nsew signal output
rlabel metal2 s 150066 -424 150122 56 8 gpio_analog_en[38]
port 120 nsew signal output
rlabel metal2 s 258666 -424 258722 56 8 gpio_analog_en[39]
port 121 nsew signal output
rlabel metal3 s 633270 199059 633750 199129 6 gpio_analog_en[3]
port 122 nsew signal output
rlabel metal2 s 313466 -424 313522 56 8 gpio_analog_en[40]
port 123 nsew signal output
rlabel metal2 s 368266 -424 368322 56 8 gpio_analog_en[41]
port 124 nsew signal output
rlabel metal2 s 423066 -424 423122 56 8 gpio_analog_en[42]
port 125 nsew signal output
rlabel metal2 s 477866 -424 477922 56 8 gpio_analog_en[43]
port 126 nsew signal output
rlabel metal3 s 633270 244059 633750 244129 6 gpio_analog_en[4]
port 127 nsew signal output
rlabel metal3 s 633270 289059 633750 289129 6 gpio_analog_en[5]
port 128 nsew signal output
rlabel metal3 s 633270 334259 633750 334329 6 gpio_analog_en[6]
port 129 nsew signal output
rlabel metal3 s 633270 511459 633750 511529 6 gpio_analog_en[7]
port 130 nsew signal output
rlabel metal3 s 633270 556659 633750 556729 6 gpio_analog_en[8]
port 131 nsew signal output
rlabel metal3 s 633270 601659 633750 601729 6 gpio_analog_en[9]
port 132 nsew signal output
rlabel metal3 s 633270 64947 633750 65017 6 gpio_analog_pol[0]
port 133 nsew signal output
rlabel metal3 s 633270 648147 633750 648217 6 gpio_analog_pol[10]
port 134 nsew signal output
rlabel metal3 s 633270 693147 633750 693217 6 gpio_analog_pol[11]
port 135 nsew signal output
rlabel metal3 s 633270 738147 633750 738217 6 gpio_analog_pol[12]
port 136 nsew signal output
rlabel metal3 s 633270 827347 633750 827417 6 gpio_analog_pol[13]
port 137 nsew signal output
rlabel metal3 s 633270 916547 633750 916617 6 gpio_analog_pol[14]
port 138 nsew signal output
rlabel metal2 s 592716 953270 592772 953750 6 gpio_analog_pol[15]
port 139 nsew signal output
rlabel metal2 s 490916 953270 490972 953750 6 gpio_analog_pol[16]
port 140 nsew signal output
rlabel metal2 s 439516 953270 439572 953750 6 gpio_analog_pol[17]
port 141 nsew signal output
rlabel metal2 s 350516 953270 350572 953750 6 gpio_analog_pol[18]
port 142 nsew signal output
rlabel metal2 s 248716 953270 248772 953750 6 gpio_analog_pol[19]
port 143 nsew signal output
rlabel metal3 s 633270 110147 633750 110217 6 gpio_analog_pol[1]
port 144 nsew signal output
rlabel metal2 s 197116 953270 197172 953750 6 gpio_analog_pol[20]
port 145 nsew signal output
rlabel metal2 s 145716 953270 145772 953750 6 gpio_analog_pol[21]
port 146 nsew signal output
rlabel metal2 s 94316 953270 94372 953750 6 gpio_analog_pol[22]
port 147 nsew signal output
rlabel metal2 s 42916 953270 42972 953750 6 gpio_analog_pol[23]
port 148 nsew signal output
rlabel metal3 s -424 920909 56 920979 4 gpio_analog_pol[24]
port 149 nsew signal output
rlabel metal3 s -424 751109 56 751179 4 gpio_analog_pol[25]
port 150 nsew signal output
rlabel metal3 s -424 707909 56 707979 4 gpio_analog_pol[26]
port 151 nsew signal output
rlabel metal3 s -424 664709 56 664779 4 gpio_analog_pol[27]
port 152 nsew signal output
rlabel metal3 s -424 621509 56 621579 4 gpio_analog_pol[28]
port 153 nsew signal output
rlabel metal3 s -424 578309 56 578379 4 gpio_analog_pol[29]
port 154 nsew signal output
rlabel metal3 s 633270 155147 633750 155217 6 gpio_analog_pol[2]
port 155 nsew signal output
rlabel metal3 s -424 535109 56 535179 4 gpio_analog_pol[30]
port 156 nsew signal output
rlabel metal3 s -424 491909 56 491979 4 gpio_analog_pol[31]
port 157 nsew signal output
rlabel metal3 s -424 364309 56 364379 4 gpio_analog_pol[32]
port 158 nsew signal output
rlabel metal3 s -424 321109 56 321179 4 gpio_analog_pol[33]
port 159 nsew signal output
rlabel metal3 s -424 277909 56 277979 4 gpio_analog_pol[34]
port 160 nsew signal output
rlabel metal3 s -424 234709 56 234779 4 gpio_analog_pol[35]
port 161 nsew signal output
rlabel metal3 s -424 191508 56 191580 4 gpio_analog_pol[36]
port 162 nsew signal output
rlabel metal3 s -424 148308 56 148380 4 gpio_analog_pol[37]
port 163 nsew signal output
rlabel metal2 s 151354 -424 151410 56 8 gpio_analog_pol[38]
port 164 nsew signal output
rlabel metal2 s 259954 -424 260010 56 8 gpio_analog_pol[39]
port 165 nsew signal output
rlabel metal3 s 633270 200347 633750 200417 6 gpio_analog_pol[3]
port 166 nsew signal output
rlabel metal2 s 314754 -424 314810 56 8 gpio_analog_pol[40]
port 167 nsew signal output
rlabel metal2 s 369554 -424 369610 56 8 gpio_analog_pol[41]
port 168 nsew signal output
rlabel metal2 s 424354 -424 424410 56 8 gpio_analog_pol[42]
port 169 nsew signal output
rlabel metal2 s 479154 -424 479210 56 8 gpio_analog_pol[43]
port 170 nsew signal output
rlabel metal3 s 633270 245347 633750 245417 6 gpio_analog_pol[4]
port 171 nsew signal output
rlabel metal3 s 633270 290347 633750 290417 6 gpio_analog_pol[5]
port 172 nsew signal output
rlabel metal3 s 633270 335547 633750 335617 6 gpio_analog_pol[6]
port 173 nsew signal output
rlabel metal3 s 633270 512747 633750 512817 6 gpio_analog_pol[7]
port 174 nsew signal output
rlabel metal3 s 633270 557947 633750 558017 6 gpio_analog_pol[8]
port 175 nsew signal output
rlabel metal3 s 633270 602947 633750 603017 6 gpio_analog_pol[9]
port 176 nsew signal output
rlabel metal3 s 633270 67983 633750 68053 6 gpio_analog_sel[0]
port 177 nsew signal output
rlabel metal3 s 633270 651183 633750 651253 6 gpio_analog_sel[10]
port 178 nsew signal output
rlabel metal3 s 633270 696183 633750 696253 6 gpio_analog_sel[11]
port 179 nsew signal output
rlabel metal3 s 633270 741183 633750 741253 6 gpio_analog_sel[12]
port 180 nsew signal output
rlabel metal3 s 633270 830383 633750 830453 6 gpio_analog_sel[13]
port 181 nsew signal output
rlabel metal3 s 633270 919583 633750 919653 6 gpio_analog_sel[14]
port 182 nsew signal output
rlabel metal2 s 589680 953270 589736 953750 6 gpio_analog_sel[15]
port 183 nsew signal output
rlabel metal2 s 487880 953270 487936 953750 6 gpio_analog_sel[16]
port 184 nsew signal output
rlabel metal2 s 436480 953270 436536 953750 6 gpio_analog_sel[17]
port 185 nsew signal output
rlabel metal2 s 347480 953270 347536 953750 6 gpio_analog_sel[18]
port 186 nsew signal output
rlabel metal2 s 245680 953270 245736 953750 6 gpio_analog_sel[19]
port 187 nsew signal output
rlabel metal3 s 633270 113183 633750 113253 6 gpio_analog_sel[1]
port 188 nsew signal output
rlabel metal2 s 194080 953270 194136 953750 6 gpio_analog_sel[20]
port 189 nsew signal output
rlabel metal2 s 142680 953270 142736 953750 6 gpio_analog_sel[21]
port 190 nsew signal output
rlabel metal2 s 91280 953270 91336 953750 6 gpio_analog_sel[22]
port 191 nsew signal output
rlabel metal2 s 39880 953270 39936 953750 6 gpio_analog_sel[23]
port 192 nsew signal output
rlabel metal3 s -424 917873 56 917943 4 gpio_analog_sel[24]
port 193 nsew signal output
rlabel metal3 s -424 748073 56 748143 4 gpio_analog_sel[25]
port 194 nsew signal output
rlabel metal3 s -424 704873 56 704943 4 gpio_analog_sel[26]
port 195 nsew signal output
rlabel metal3 s -424 661673 56 661743 4 gpio_analog_sel[27]
port 196 nsew signal output
rlabel metal3 s -424 618473 56 618543 4 gpio_analog_sel[28]
port 197 nsew signal output
rlabel metal3 s -424 575273 56 575343 4 gpio_analog_sel[29]
port 198 nsew signal output
rlabel metal3 s 633270 158183 633750 158253 6 gpio_analog_sel[2]
port 199 nsew signal output
rlabel metal3 s -424 532073 56 532143 4 gpio_analog_sel[30]
port 200 nsew signal output
rlabel metal3 s -424 488873 56 488943 4 gpio_analog_sel[31]
port 201 nsew signal output
rlabel metal3 s -424 361273 56 361343 4 gpio_analog_sel[32]
port 202 nsew signal output
rlabel metal3 s -424 318073 56 318143 4 gpio_analog_sel[33]
port 203 nsew signal output
rlabel metal3 s -424 274873 56 274943 4 gpio_analog_sel[34]
port 204 nsew signal output
rlabel metal3 s -424 231673 56 231743 4 gpio_analog_sel[35]
port 205 nsew signal output
rlabel metal3 s -424 188472 56 188544 4 gpio_analog_sel[36]
port 206 nsew signal output
rlabel metal3 s -424 145272 56 145344 4 gpio_analog_sel[37]
port 207 nsew signal output
rlabel metal2 s 154390 -424 154446 56 8 gpio_analog_sel[38]
port 208 nsew signal output
rlabel metal2 s 262990 -424 263046 56 8 gpio_analog_sel[39]
port 209 nsew signal output
rlabel metal3 s 633270 203383 633750 203453 6 gpio_analog_sel[3]
port 210 nsew signal output
rlabel metal2 s 317790 -424 317846 56 8 gpio_analog_sel[40]
port 211 nsew signal output
rlabel metal2 s 372590 -424 372646 56 8 gpio_analog_sel[41]
port 212 nsew signal output
rlabel metal2 s 427390 -424 427446 56 8 gpio_analog_sel[42]
port 213 nsew signal output
rlabel metal2 s 482190 -424 482246 56 8 gpio_analog_sel[43]
port 214 nsew signal output
rlabel metal3 s 633270 248383 633750 248453 6 gpio_analog_sel[4]
port 215 nsew signal output
rlabel metal3 s 633270 293383 633750 293453 6 gpio_analog_sel[5]
port 216 nsew signal output
rlabel metal3 s 633270 338583 633750 338653 6 gpio_analog_sel[6]
port 217 nsew signal output
rlabel metal3 s 633270 515783 633750 515853 6 gpio_analog_sel[7]
port 218 nsew signal output
rlabel metal3 s 633270 560983 633750 561053 6 gpio_analog_sel[8]
port 219 nsew signal output
rlabel metal3 s 633270 605983 633750 606053 6 gpio_analog_sel[9]
port 220 nsew signal output
rlabel metal3 s 633270 64303 633750 64373 6 gpio_dm0[0]
port 221 nsew signal output
rlabel metal3 s 633270 647503 633750 647573 6 gpio_dm0[10]
port 222 nsew signal output
rlabel metal3 s 633270 692503 633750 692573 6 gpio_dm0[11]
port 223 nsew signal output
rlabel metal3 s 633270 737503 633750 737573 6 gpio_dm0[12]
port 224 nsew signal output
rlabel metal3 s 633270 826703 633750 826773 6 gpio_dm0[13]
port 225 nsew signal output
rlabel metal3 s 633270 915903 633750 915973 6 gpio_dm0[14]
port 226 nsew signal output
rlabel metal2 s 593360 953270 593416 953750 6 gpio_dm0[15]
port 227 nsew signal output
rlabel metal2 s 491560 953270 491616 953750 6 gpio_dm0[16]
port 228 nsew signal output
rlabel metal2 s 440160 953270 440216 953750 6 gpio_dm0[17]
port 229 nsew signal output
rlabel metal2 s 351160 953270 351216 953750 6 gpio_dm0[18]
port 230 nsew signal output
rlabel metal2 s 249360 953270 249416 953750 6 gpio_dm0[19]
port 231 nsew signal output
rlabel metal3 s 633270 109503 633750 109573 6 gpio_dm0[1]
port 232 nsew signal output
rlabel metal2 s 197760 953270 197816 953750 6 gpio_dm0[20]
port 233 nsew signal output
rlabel metal2 s 146360 953270 146416 953750 6 gpio_dm0[21]
port 234 nsew signal output
rlabel metal2 s 94960 953270 95016 953750 6 gpio_dm0[22]
port 235 nsew signal output
rlabel metal2 s 43560 953270 43616 953750 6 gpio_dm0[23]
port 236 nsew signal output
rlabel metal3 s -424 921553 56 921623 4 gpio_dm0[24]
port 237 nsew signal output
rlabel metal3 s -424 751753 56 751823 4 gpio_dm0[25]
port 238 nsew signal output
rlabel metal3 s -424 708553 56 708623 4 gpio_dm0[26]
port 239 nsew signal output
rlabel metal3 s -424 665353 56 665423 4 gpio_dm0[27]
port 240 nsew signal output
rlabel metal3 s -424 622153 56 622223 4 gpio_dm0[28]
port 241 nsew signal output
rlabel metal3 s -424 578953 56 579023 4 gpio_dm0[29]
port 242 nsew signal output
rlabel metal3 s 633270 154503 633750 154573 6 gpio_dm0[2]
port 243 nsew signal output
rlabel metal3 s -424 535753 56 535823 4 gpio_dm0[30]
port 244 nsew signal output
rlabel metal3 s -424 492553 56 492623 4 gpio_dm0[31]
port 245 nsew signal output
rlabel metal3 s -424 364953 56 365023 4 gpio_dm0[32]
port 246 nsew signal output
rlabel metal3 s -424 321753 56 321823 4 gpio_dm0[33]
port 247 nsew signal output
rlabel metal3 s -424 278553 56 278623 4 gpio_dm0[34]
port 248 nsew signal output
rlabel metal3 s -424 235353 56 235423 4 gpio_dm0[35]
port 249 nsew signal output
rlabel metal3 s -424 192152 56 192224 4 gpio_dm0[36]
port 250 nsew signal output
rlabel metal3 s -424 148952 56 149024 4 gpio_dm0[37]
port 251 nsew signal output
rlabel metal2 s 148870 -424 148926 56 8 gpio_dm0[38]
port 252 nsew signal output
rlabel metal2 s 259310 -424 259366 56 8 gpio_dm0[39]
port 253 nsew signal output
rlabel metal3 s 633270 199703 633750 199773 6 gpio_dm0[3]
port 254 nsew signal output
rlabel metal2 s 314110 -424 314166 56 8 gpio_dm0[40]
port 255 nsew signal output
rlabel metal2 s 368910 -424 368966 56 8 gpio_dm0[41]
port 256 nsew signal output
rlabel metal2 s 423710 -424 423766 56 8 gpio_dm0[42]
port 257 nsew signal output
rlabel metal2 s 478510 -424 478566 56 8 gpio_dm0[43]
port 258 nsew signal output
rlabel metal3 s 633270 244703 633750 244773 6 gpio_dm0[4]
port 259 nsew signal output
rlabel metal3 s 633270 289703 633750 289773 6 gpio_dm0[5]
port 260 nsew signal output
rlabel metal3 s 633270 334903 633750 334973 6 gpio_dm0[6]
port 261 nsew signal output
rlabel metal3 s 633270 512103 633750 512173 6 gpio_dm0[7]
port 262 nsew signal output
rlabel metal3 s 633270 557303 633750 557373 6 gpio_dm0[8]
port 263 nsew signal output
rlabel metal3 s 633270 602303 633750 602373 6 gpio_dm0[9]
port 264 nsew signal output
rlabel metal3 s 633270 62463 633750 62533 6 gpio_dm1[0]
port 265 nsew signal output
rlabel metal3 s 633270 645663 633750 645733 6 gpio_dm1[10]
port 266 nsew signal output
rlabel metal3 s 633270 690663 633750 690733 6 gpio_dm1[11]
port 267 nsew signal output
rlabel metal3 s 633270 735663 633750 735733 6 gpio_dm1[12]
port 268 nsew signal output
rlabel metal3 s 633270 824863 633750 824933 6 gpio_dm1[13]
port 269 nsew signal output
rlabel metal3 s 633270 914063 633750 914133 6 gpio_dm1[14]
port 270 nsew signal output
rlabel metal2 s 595200 953270 595256 953750 6 gpio_dm1[15]
port 271 nsew signal output
rlabel metal2 s 493400 953270 493456 953750 6 gpio_dm1[16]
port 272 nsew signal output
rlabel metal2 s 442000 953270 442056 953750 6 gpio_dm1[17]
port 273 nsew signal output
rlabel metal2 s 353000 953270 353056 953750 6 gpio_dm1[18]
port 274 nsew signal output
rlabel metal2 s 251200 953270 251256 953750 6 gpio_dm1[19]
port 275 nsew signal output
rlabel metal3 s 633270 107663 633750 107733 6 gpio_dm1[1]
port 276 nsew signal output
rlabel metal2 s 199600 953270 199656 953750 6 gpio_dm1[20]
port 277 nsew signal output
rlabel metal2 s 148200 953270 148256 953750 6 gpio_dm1[21]
port 278 nsew signal output
rlabel metal2 s 96800 953270 96856 953750 6 gpio_dm1[22]
port 279 nsew signal output
rlabel metal2 s 45400 953270 45456 953750 6 gpio_dm1[23]
port 280 nsew signal output
rlabel metal3 s -424 923393 56 923463 4 gpio_dm1[24]
port 281 nsew signal output
rlabel metal3 s -424 753593 56 753663 4 gpio_dm1[25]
port 282 nsew signal output
rlabel metal3 s -424 710393 56 710463 4 gpio_dm1[26]
port 283 nsew signal output
rlabel metal3 s -424 667193 56 667263 4 gpio_dm1[27]
port 284 nsew signal output
rlabel metal3 s -424 623993 56 624063 4 gpio_dm1[28]
port 285 nsew signal output
rlabel metal3 s -424 580793 56 580863 4 gpio_dm1[29]
port 286 nsew signal output
rlabel metal3 s 633270 152663 633750 152733 6 gpio_dm1[2]
port 287 nsew signal output
rlabel metal3 s -424 537593 56 537663 4 gpio_dm1[30]
port 288 nsew signal output
rlabel metal3 s -424 494393 56 494463 4 gpio_dm1[31]
port 289 nsew signal output
rlabel metal3 s -424 366793 56 366863 4 gpio_dm1[32]
port 290 nsew signal output
rlabel metal3 s -424 323593 56 323663 4 gpio_dm1[33]
port 291 nsew signal output
rlabel metal3 s -424 280393 56 280463 4 gpio_dm1[34]
port 292 nsew signal output
rlabel metal3 s -424 237193 56 237263 4 gpio_dm1[35]
port 293 nsew signal output
rlabel metal3 s -424 193992 56 194064 4 gpio_dm1[36]
port 294 nsew signal output
rlabel metal3 s -424 150792 56 150864 4 gpio_dm1[37]
port 295 nsew signal output
rlabel metal2 s 150710 -424 150766 56 8 gpio_dm1[38]
port 296 nsew signal output
rlabel metal2 s 257470 -424 257526 56 8 gpio_dm1[39]
port 297 nsew signal output
rlabel metal3 s 633270 197863 633750 197933 6 gpio_dm1[3]
port 298 nsew signal output
rlabel metal2 s 312270 -424 312326 56 8 gpio_dm1[40]
port 299 nsew signal output
rlabel metal2 s 367070 -424 367126 56 8 gpio_dm1[41]
port 300 nsew signal output
rlabel metal2 s 421870 -424 421926 56 8 gpio_dm1[42]
port 301 nsew signal output
rlabel metal2 s 476670 -424 476726 56 8 gpio_dm1[43]
port 302 nsew signal output
rlabel metal3 s 633270 242863 633750 242933 6 gpio_dm1[4]
port 303 nsew signal output
rlabel metal3 s 633270 287863 633750 287933 6 gpio_dm1[5]
port 304 nsew signal output
rlabel metal3 s 633270 333063 633750 333133 6 gpio_dm1[6]
port 305 nsew signal output
rlabel metal3 s 633270 510263 633750 510333 6 gpio_dm1[7]
port 306 nsew signal output
rlabel metal3 s 633270 555463 633750 555533 6 gpio_dm1[8]
port 307 nsew signal output
rlabel metal3 s 633270 600463 633750 600533 6 gpio_dm1[9]
port 308 nsew signal output
rlabel metal3 s 633270 68627 633750 68697 6 gpio_dm2[0]
port 309 nsew signal output
rlabel metal3 s 633270 651827 633750 651897 6 gpio_dm2[10]
port 310 nsew signal output
rlabel metal3 s 633270 696827 633750 696897 6 gpio_dm2[11]
port 311 nsew signal output
rlabel metal3 s 633270 741827 633750 741897 6 gpio_dm2[12]
port 312 nsew signal output
rlabel metal3 s 633270 831027 633750 831097 6 gpio_dm2[13]
port 313 nsew signal output
rlabel metal3 s 633270 920227 633750 920297 6 gpio_dm2[14]
port 314 nsew signal output
rlabel metal2 s 589036 953270 589092 953750 6 gpio_dm2[15]
port 315 nsew signal output
rlabel metal2 s 487236 953270 487292 953750 6 gpio_dm2[16]
port 316 nsew signal output
rlabel metal2 s 435836 953270 435892 953750 6 gpio_dm2[17]
port 317 nsew signal output
rlabel metal2 s 346836 953270 346892 953750 6 gpio_dm2[18]
port 318 nsew signal output
rlabel metal2 s 245036 953270 245092 953750 6 gpio_dm2[19]
port 319 nsew signal output
rlabel metal3 s 633270 113827 633750 113897 6 gpio_dm2[1]
port 320 nsew signal output
rlabel metal2 s 193436 953270 193492 953750 6 gpio_dm2[20]
port 321 nsew signal output
rlabel metal2 s 142036 953270 142092 953750 6 gpio_dm2[21]
port 322 nsew signal output
rlabel metal2 s 90636 953270 90692 953750 6 gpio_dm2[22]
port 323 nsew signal output
rlabel metal2 s 39236 953270 39292 953750 6 gpio_dm2[23]
port 324 nsew signal output
rlabel metal3 s -424 917229 56 917299 4 gpio_dm2[24]
port 325 nsew signal output
rlabel metal3 s -424 747429 56 747499 4 gpio_dm2[25]
port 326 nsew signal output
rlabel metal3 s -424 704229 56 704299 4 gpio_dm2[26]
port 327 nsew signal output
rlabel metal3 s -424 661029 56 661099 4 gpio_dm2[27]
port 328 nsew signal output
rlabel metal3 s -424 617829 56 617899 4 gpio_dm2[28]
port 329 nsew signal output
rlabel metal3 s -424 574629 56 574699 4 gpio_dm2[29]
port 330 nsew signal output
rlabel metal3 s 633270 158827 633750 158897 6 gpio_dm2[2]
port 331 nsew signal output
rlabel metal3 s -424 531429 56 531499 4 gpio_dm2[30]
port 332 nsew signal output
rlabel metal3 s -424 488229 56 488299 4 gpio_dm2[31]
port 333 nsew signal output
rlabel metal3 s -424 360629 56 360699 4 gpio_dm2[32]
port 334 nsew signal output
rlabel metal3 s -424 317429 56 317499 4 gpio_dm2[33]
port 335 nsew signal output
rlabel metal3 s -424 274229 56 274299 4 gpio_dm2[34]
port 336 nsew signal output
rlabel metal3 s -424 231029 56 231099 4 gpio_dm2[35]
port 337 nsew signal output
rlabel metal3 s -424 187828 56 187900 4 gpio_dm2[36]
port 338 nsew signal output
rlabel metal3 s -424 144628 56 144700 4 gpio_dm2[37]
port 339 nsew signal output
rlabel metal2 s 155034 -424 155090 56 8 gpio_dm2[38]
port 340 nsew signal output
rlabel metal2 s 263634 -424 263690 56 8 gpio_dm2[39]
port 341 nsew signal output
rlabel metal3 s 633270 204027 633750 204097 6 gpio_dm2[3]
port 342 nsew signal output
rlabel metal2 s 318434 -424 318490 56 8 gpio_dm2[40]
port 343 nsew signal output
rlabel metal2 s 373234 -424 373290 56 8 gpio_dm2[41]
port 344 nsew signal output
rlabel metal2 s 428034 -424 428090 56 8 gpio_dm2[42]
port 345 nsew signal output
rlabel metal2 s 482834 -424 482890 56 8 gpio_dm2[43]
port 346 nsew signal output
rlabel metal3 s 633270 249027 633750 249097 6 gpio_dm2[4]
port 347 nsew signal output
rlabel metal3 s 633270 294027 633750 294097 6 gpio_dm2[5]
port 348 nsew signal output
rlabel metal3 s 633270 339227 633750 339297 6 gpio_dm2[6]
port 349 nsew signal output
rlabel metal3 s 633270 516427 633750 516497 6 gpio_dm2[7]
port 350 nsew signal output
rlabel metal3 s 633270 561627 633750 561697 6 gpio_dm2[8]
port 351 nsew signal output
rlabel metal3 s 633270 606627 633750 606697 6 gpio_dm2[9]
port 352 nsew signal output
rlabel metal3 s 633270 69271 633750 69341 6 gpio_holdover[0]
port 353 nsew signal output
rlabel metal3 s 633270 652471 633750 652541 6 gpio_holdover[10]
port 354 nsew signal output
rlabel metal3 s 633270 697471 633750 697541 6 gpio_holdover[11]
port 355 nsew signal output
rlabel metal3 s 633270 742471 633750 742541 6 gpio_holdover[12]
port 356 nsew signal output
rlabel metal3 s 633270 831671 633750 831741 6 gpio_holdover[13]
port 357 nsew signal output
rlabel metal3 s 633270 920871 633750 920941 6 gpio_holdover[14]
port 358 nsew signal output
rlabel metal2 s 588392 953270 588448 953750 6 gpio_holdover[15]
port 359 nsew signal output
rlabel metal2 s 486592 953270 486648 953750 6 gpio_holdover[16]
port 360 nsew signal output
rlabel metal2 s 435192 953270 435248 953750 6 gpio_holdover[17]
port 361 nsew signal output
rlabel metal2 s 346192 953270 346248 953750 6 gpio_holdover[18]
port 362 nsew signal output
rlabel metal2 s 244392 953270 244448 953750 6 gpio_holdover[19]
port 363 nsew signal output
rlabel metal3 s 633270 114471 633750 114541 6 gpio_holdover[1]
port 364 nsew signal output
rlabel metal2 s 192792 953270 192848 953750 6 gpio_holdover[20]
port 365 nsew signal output
rlabel metal2 s 141392 953270 141448 953750 6 gpio_holdover[21]
port 366 nsew signal output
rlabel metal2 s 89992 953270 90048 953750 6 gpio_holdover[22]
port 367 nsew signal output
rlabel metal2 s 38592 953270 38648 953750 6 gpio_holdover[23]
port 368 nsew signal output
rlabel metal3 s -424 916585 56 916655 4 gpio_holdover[24]
port 369 nsew signal output
rlabel metal3 s -424 746785 56 746855 4 gpio_holdover[25]
port 370 nsew signal output
rlabel metal3 s -424 703585 56 703655 4 gpio_holdover[26]
port 371 nsew signal output
rlabel metal3 s -424 660385 56 660455 4 gpio_holdover[27]
port 372 nsew signal output
rlabel metal3 s -424 617185 56 617255 4 gpio_holdover[28]
port 373 nsew signal output
rlabel metal3 s -424 573985 56 574055 4 gpio_holdover[29]
port 374 nsew signal output
rlabel metal3 s 633270 159471 633750 159541 6 gpio_holdover[2]
port 375 nsew signal output
rlabel metal3 s -424 530785 56 530855 4 gpio_holdover[30]
port 376 nsew signal output
rlabel metal3 s -424 487585 56 487655 4 gpio_holdover[31]
port 377 nsew signal output
rlabel metal3 s -424 359985 56 360055 4 gpio_holdover[32]
port 378 nsew signal output
rlabel metal3 s -424 316785 56 316855 4 gpio_holdover[33]
port 379 nsew signal output
rlabel metal3 s -424 273585 56 273655 4 gpio_holdover[34]
port 380 nsew signal output
rlabel metal3 s -424 230385 56 230455 4 gpio_holdover[35]
port 381 nsew signal output
rlabel metal3 s -424 187184 56 187256 4 gpio_holdover[36]
port 382 nsew signal output
rlabel metal3 s -424 143984 56 144056 4 gpio_holdover[37]
port 383 nsew signal output
rlabel metal2 s 155678 -424 155734 56 8 gpio_holdover[38]
port 384 nsew signal output
rlabel metal2 s 264278 -424 264334 56 8 gpio_holdover[39]
port 385 nsew signal output
rlabel metal3 s 633270 204671 633750 204741 6 gpio_holdover[3]
port 386 nsew signal output
rlabel metal2 s 319078 -424 319134 56 8 gpio_holdover[40]
port 387 nsew signal output
rlabel metal2 s 373878 -424 373934 56 8 gpio_holdover[41]
port 388 nsew signal output
rlabel metal2 s 428678 -424 428734 56 8 gpio_holdover[42]
port 389 nsew signal output
rlabel metal2 s 483478 -424 483534 56 8 gpio_holdover[43]
port 390 nsew signal output
rlabel metal3 s 633270 249671 633750 249741 6 gpio_holdover[4]
port 391 nsew signal output
rlabel metal3 s 633270 294671 633750 294741 6 gpio_holdover[5]
port 392 nsew signal output
rlabel metal3 s 633270 339871 633750 339941 6 gpio_holdover[6]
port 393 nsew signal output
rlabel metal3 s 633270 517071 633750 517141 6 gpio_holdover[7]
port 394 nsew signal output
rlabel metal3 s 633270 562271 633750 562341 6 gpio_holdover[8]
port 395 nsew signal output
rlabel metal3 s 633270 607271 633750 607341 6 gpio_holdover[9]
port 396 nsew signal output
rlabel metal3 s 633270 72307 633750 72377 6 gpio_ib_mode_sel[0]
port 397 nsew signal output
rlabel metal3 s 633270 655507 633750 655577 6 gpio_ib_mode_sel[10]
port 398 nsew signal output
rlabel metal3 s 633270 700507 633750 700577 6 gpio_ib_mode_sel[11]
port 399 nsew signal output
rlabel metal3 s 633270 745507 633750 745577 6 gpio_ib_mode_sel[12]
port 400 nsew signal output
rlabel metal3 s 633270 834707 633750 834777 6 gpio_ib_mode_sel[13]
port 401 nsew signal output
rlabel metal3 s 633270 923907 633750 923977 6 gpio_ib_mode_sel[14]
port 402 nsew signal output
rlabel metal2 s 585356 953270 585412 953750 6 gpio_ib_mode_sel[15]
port 403 nsew signal output
rlabel metal2 s 483556 953270 483612 953750 6 gpio_ib_mode_sel[16]
port 404 nsew signal output
rlabel metal2 s 432156 953270 432212 953750 6 gpio_ib_mode_sel[17]
port 405 nsew signal output
rlabel metal2 s 343156 953270 343212 953750 6 gpio_ib_mode_sel[18]
port 406 nsew signal output
rlabel metal2 s 241356 953270 241412 953750 6 gpio_ib_mode_sel[19]
port 407 nsew signal output
rlabel metal3 s 633270 117507 633750 117577 6 gpio_ib_mode_sel[1]
port 408 nsew signal output
rlabel metal2 s 189756 953270 189812 953750 6 gpio_ib_mode_sel[20]
port 409 nsew signal output
rlabel metal2 s 138356 953270 138412 953750 6 gpio_ib_mode_sel[21]
port 410 nsew signal output
rlabel metal2 s 86956 953270 87012 953750 6 gpio_ib_mode_sel[22]
port 411 nsew signal output
rlabel metal2 s 35556 953270 35612 953750 6 gpio_ib_mode_sel[23]
port 412 nsew signal output
rlabel metal3 s -424 913549 56 913619 4 gpio_ib_mode_sel[24]
port 413 nsew signal output
rlabel metal3 s -424 743749 56 743819 4 gpio_ib_mode_sel[25]
port 414 nsew signal output
rlabel metal3 s -424 700549 56 700619 4 gpio_ib_mode_sel[26]
port 415 nsew signal output
rlabel metal3 s -424 657349 56 657419 4 gpio_ib_mode_sel[27]
port 416 nsew signal output
rlabel metal3 s -424 614149 56 614219 4 gpio_ib_mode_sel[28]
port 417 nsew signal output
rlabel metal3 s -424 570949 56 571019 4 gpio_ib_mode_sel[29]
port 418 nsew signal output
rlabel metal3 s 633270 162507 633750 162577 6 gpio_ib_mode_sel[2]
port 419 nsew signal output
rlabel metal3 s -424 527749 56 527819 4 gpio_ib_mode_sel[30]
port 420 nsew signal output
rlabel metal3 s -424 484549 56 484619 4 gpio_ib_mode_sel[31]
port 421 nsew signal output
rlabel metal3 s -424 356949 56 357019 4 gpio_ib_mode_sel[32]
port 422 nsew signal output
rlabel metal3 s -424 313749 56 313819 4 gpio_ib_mode_sel[33]
port 423 nsew signal output
rlabel metal3 s -424 270549 56 270619 4 gpio_ib_mode_sel[34]
port 424 nsew signal output
rlabel metal3 s -424 227349 56 227419 4 gpio_ib_mode_sel[35]
port 425 nsew signal output
rlabel metal3 s -424 184148 56 184220 4 gpio_ib_mode_sel[36]
port 426 nsew signal output
rlabel metal3 s -424 140948 56 141020 4 gpio_ib_mode_sel[37]
port 427 nsew signal output
rlabel metal2 s 158714 -424 158770 56 8 gpio_ib_mode_sel[38]
port 428 nsew signal output
rlabel metal2 s 267314 -424 267370 56 8 gpio_ib_mode_sel[39]
port 429 nsew signal output
rlabel metal3 s 633270 207707 633750 207777 6 gpio_ib_mode_sel[3]
port 430 nsew signal output
rlabel metal2 s 322114 -424 322170 56 8 gpio_ib_mode_sel[40]
port 431 nsew signal output
rlabel metal2 s 376914 -424 376970 56 8 gpio_ib_mode_sel[41]
port 432 nsew signal output
rlabel metal2 s 431714 -424 431770 56 8 gpio_ib_mode_sel[42]
port 433 nsew signal output
rlabel metal2 s 486514 -424 486570 56 8 gpio_ib_mode_sel[43]
port 434 nsew signal output
rlabel metal3 s 633270 252707 633750 252777 6 gpio_ib_mode_sel[4]
port 435 nsew signal output
rlabel metal3 s 633270 297707 633750 297777 6 gpio_ib_mode_sel[5]
port 436 nsew signal output
rlabel metal3 s 633270 342907 633750 342977 6 gpio_ib_mode_sel[6]
port 437 nsew signal output
rlabel metal3 s 633270 520107 633750 520177 6 gpio_ib_mode_sel[7]
port 438 nsew signal output
rlabel metal3 s 633270 565307 633750 565377 6 gpio_ib_mode_sel[8]
port 439 nsew signal output
rlabel metal3 s 633270 610307 633750 610377 6 gpio_ib_mode_sel[9]
port 440 nsew signal output
rlabel metal3 s 633270 58783 633750 58853 6 gpio_in[0]
port 441 nsew signal input
rlabel metal3 s 633270 641983 633750 642053 6 gpio_in[10]
port 442 nsew signal input
rlabel metal3 s 633270 686983 633750 687053 6 gpio_in[11]
port 443 nsew signal input
rlabel metal3 s 633270 731983 633750 732053 6 gpio_in[12]
port 444 nsew signal input
rlabel metal3 s 633270 821183 633750 821253 6 gpio_in[13]
port 445 nsew signal input
rlabel metal3 s 633270 910383 633750 910453 6 gpio_in[14]
port 446 nsew signal input
rlabel metal2 s 598880 953270 598936 953750 6 gpio_in[15]
port 447 nsew signal input
rlabel metal2 s 497080 953270 497136 953750 6 gpio_in[16]
port 448 nsew signal input
rlabel metal2 s 445680 953270 445736 953750 6 gpio_in[17]
port 449 nsew signal input
rlabel metal2 s 356680 953270 356736 953750 6 gpio_in[18]
port 450 nsew signal input
rlabel metal2 s 254880 953270 254936 953750 6 gpio_in[19]
port 451 nsew signal input
rlabel metal3 s 633270 103983 633750 104053 6 gpio_in[1]
port 452 nsew signal input
rlabel metal2 s 203280 953270 203336 953750 6 gpio_in[20]
port 453 nsew signal input
rlabel metal2 s 151880 953270 151936 953750 6 gpio_in[21]
port 454 nsew signal input
rlabel metal2 s 100480 953270 100536 953750 6 gpio_in[22]
port 455 nsew signal input
rlabel metal2 s 49080 953270 49136 953750 6 gpio_in[23]
port 456 nsew signal input
rlabel metal3 s -424 927073 56 927143 4 gpio_in[24]
port 457 nsew signal input
rlabel metal3 s -424 757273 56 757343 4 gpio_in[25]
port 458 nsew signal input
rlabel metal3 s -424 714073 56 714143 4 gpio_in[26]
port 459 nsew signal input
rlabel metal3 s -424 670873 56 670943 4 gpio_in[27]
port 460 nsew signal input
rlabel metal3 s -424 627673 56 627743 4 gpio_in[28]
port 461 nsew signal input
rlabel metal3 s -424 584473 56 584543 4 gpio_in[29]
port 462 nsew signal input
rlabel metal3 s 633270 148983 633750 149053 6 gpio_in[2]
port 463 nsew signal input
rlabel metal3 s -424 541273 56 541343 4 gpio_in[30]
port 464 nsew signal input
rlabel metal3 s -424 498073 56 498143 4 gpio_in[31]
port 465 nsew signal input
rlabel metal3 s -424 370473 56 370543 4 gpio_in[32]
port 466 nsew signal input
rlabel metal3 s -424 327273 56 327343 4 gpio_in[33]
port 467 nsew signal input
rlabel metal3 s -424 284073 56 284143 4 gpio_in[34]
port 468 nsew signal input
rlabel metal3 s -424 240873 56 240943 4 gpio_in[35]
port 469 nsew signal input
rlabel metal3 s -424 197672 56 197744 4 gpio_in[36]
port 470 nsew signal input
rlabel metal3 s -424 154472 56 154544 4 gpio_in[37]
port 471 nsew signal input
rlabel metal2 s 145190 -424 145246 56 8 gpio_in[38]
port 472 nsew signal input
rlabel metal2 s 253790 -424 253846 56 8 gpio_in[39]
port 473 nsew signal input
rlabel metal3 s 633270 194183 633750 194253 6 gpio_in[3]
port 474 nsew signal input
rlabel metal2 s 308590 -424 308646 56 8 gpio_in[40]
port 475 nsew signal input
rlabel metal2 s 363390 -424 363446 56 8 gpio_in[41]
port 476 nsew signal input
rlabel metal2 s 418190 -424 418246 56 8 gpio_in[42]
port 477 nsew signal input
rlabel metal2 s 472990 -424 473046 56 8 gpio_in[43]
port 478 nsew signal input
rlabel metal3 s 633270 239183 633750 239253 6 gpio_in[4]
port 479 nsew signal input
rlabel metal3 s 633270 284183 633750 284253 6 gpio_in[5]
port 480 nsew signal input
rlabel metal3 s 633270 329383 633750 329453 6 gpio_in[6]
port 481 nsew signal input
rlabel metal3 s 633270 506583 633750 506653 6 gpio_in[7]
port 482 nsew signal input
rlabel metal3 s 633270 551783 633750 551853 6 gpio_in[8]
port 483 nsew signal input
rlabel metal3 s 633270 596783 633750 596853 6 gpio_in[9]
port 484 nsew signal input
rlabel metal3 s 633270 73503 633750 73573 6 gpio_in_h[0]
port 485 nsew signal input
rlabel metal3 s 633270 656703 633750 656773 6 gpio_in_h[10]
port 486 nsew signal input
rlabel metal3 s 633270 701703 633750 701773 6 gpio_in_h[11]
port 487 nsew signal input
rlabel metal3 s 633270 746703 633750 746773 6 gpio_in_h[12]
port 488 nsew signal input
rlabel metal3 s 633270 835903 633750 835973 6 gpio_in_h[13]
port 489 nsew signal input
rlabel metal3 s 633270 925103 633750 925173 6 gpio_in_h[14]
port 490 nsew signal input
rlabel metal2 s 584160 953270 584216 953750 6 gpio_in_h[15]
port 491 nsew signal input
rlabel metal2 s 482360 953270 482416 953750 6 gpio_in_h[16]
port 492 nsew signal input
rlabel metal2 s 430960 953270 431016 953750 6 gpio_in_h[17]
port 493 nsew signal input
rlabel metal2 s 341960 953270 342016 953750 6 gpio_in_h[18]
port 494 nsew signal input
rlabel metal2 s 240160 953270 240216 953750 6 gpio_in_h[19]
port 495 nsew signal input
rlabel metal3 s 633270 118703 633750 118773 6 gpio_in_h[1]
port 496 nsew signal input
rlabel metal2 s 188560 953270 188616 953750 6 gpio_in_h[20]
port 497 nsew signal input
rlabel metal2 s 137160 953270 137216 953750 6 gpio_in_h[21]
port 498 nsew signal input
rlabel metal2 s 85760 953270 85816 953750 6 gpio_in_h[22]
port 499 nsew signal input
rlabel metal2 s 34360 953270 34416 953750 6 gpio_in_h[23]
port 500 nsew signal input
rlabel metal3 s -424 912353 56 912423 4 gpio_in_h[24]
port 501 nsew signal input
rlabel metal3 s -424 742553 56 742623 4 gpio_in_h[25]
port 502 nsew signal input
rlabel metal3 s -424 699353 56 699423 4 gpio_in_h[26]
port 503 nsew signal input
rlabel metal3 s -424 656153 56 656223 4 gpio_in_h[27]
port 504 nsew signal input
rlabel metal3 s -424 612953 56 613023 4 gpio_in_h[28]
port 505 nsew signal input
rlabel metal3 s -424 569753 56 569823 4 gpio_in_h[29]
port 506 nsew signal input
rlabel metal3 s 633270 163703 633750 163773 6 gpio_in_h[2]
port 507 nsew signal input
rlabel metal3 s -424 526553 56 526623 4 gpio_in_h[30]
port 508 nsew signal input
rlabel metal3 s -424 483353 56 483423 4 gpio_in_h[31]
port 509 nsew signal input
rlabel metal3 s -424 355753 56 355823 4 gpio_in_h[32]
port 510 nsew signal input
rlabel metal3 s -424 312553 56 312623 4 gpio_in_h[33]
port 511 nsew signal input
rlabel metal3 s -424 269353 56 269423 4 gpio_in_h[34]
port 512 nsew signal input
rlabel metal3 s -424 226153 56 226223 4 gpio_in_h[35]
port 513 nsew signal input
rlabel metal3 s -424 182952 56 183024 4 gpio_in_h[36]
port 514 nsew signal input
rlabel metal3 s -424 139752 56 139824 4 gpio_in_h[37]
port 515 nsew signal input
rlabel metal2 s 159910 -424 159966 56 8 gpio_in_h[38]
port 516 nsew signal input
rlabel metal2 s 268510 -424 268566 56 8 gpio_in_h[39]
port 517 nsew signal input
rlabel metal3 s 633270 208903 633750 208973 6 gpio_in_h[3]
port 518 nsew signal input
rlabel metal2 s 323310 -424 323366 56 8 gpio_in_h[40]
port 519 nsew signal input
rlabel metal2 s 378110 -424 378166 56 8 gpio_in_h[41]
port 520 nsew signal input
rlabel metal2 s 432910 -424 432966 56 8 gpio_in_h[42]
port 521 nsew signal input
rlabel metal2 s 487710 -424 487766 56 8 gpio_in_h[43]
port 522 nsew signal input
rlabel metal3 s 633270 253903 633750 253973 6 gpio_in_h[4]
port 523 nsew signal input
rlabel metal3 s 633270 298903 633750 298973 6 gpio_in_h[5]
port 524 nsew signal input
rlabel metal3 s 633270 344103 633750 344173 6 gpio_in_h[6]
port 525 nsew signal input
rlabel metal3 s 633270 521303 633750 521373 6 gpio_in_h[7]
port 526 nsew signal input
rlabel metal3 s 633270 566503 633750 566573 6 gpio_in_h[8]
port 527 nsew signal input
rlabel metal3 s 633270 611503 633750 611573 6 gpio_in_h[9]
port 528 nsew signal input
rlabel metal3 s 633270 65499 633750 65569 6 gpio_inp_dis[0]
port 529 nsew signal output
rlabel metal3 s 633270 648699 633750 648769 6 gpio_inp_dis[10]
port 530 nsew signal output
rlabel metal3 s 633270 693699 633750 693769 6 gpio_inp_dis[11]
port 531 nsew signal output
rlabel metal3 s 633270 738699 633750 738769 6 gpio_inp_dis[12]
port 532 nsew signal output
rlabel metal3 s 633270 827899 633750 827969 6 gpio_inp_dis[13]
port 533 nsew signal output
rlabel metal3 s 633270 917099 633750 917169 6 gpio_inp_dis[14]
port 534 nsew signal output
rlabel metal2 s 592164 953270 592220 953750 6 gpio_inp_dis[15]
port 535 nsew signal output
rlabel metal2 s 490364 953270 490420 953750 6 gpio_inp_dis[16]
port 536 nsew signal output
rlabel metal2 s 438964 953270 439020 953750 6 gpio_inp_dis[17]
port 537 nsew signal output
rlabel metal2 s 349964 953270 350020 953750 6 gpio_inp_dis[18]
port 538 nsew signal output
rlabel metal2 s 248164 953270 248220 953750 6 gpio_inp_dis[19]
port 539 nsew signal output
rlabel metal3 s 633270 110699 633750 110769 6 gpio_inp_dis[1]
port 540 nsew signal output
rlabel metal2 s 196564 953270 196620 953750 6 gpio_inp_dis[20]
port 541 nsew signal output
rlabel metal2 s 145164 953270 145220 953750 6 gpio_inp_dis[21]
port 542 nsew signal output
rlabel metal2 s 93764 953270 93820 953750 6 gpio_inp_dis[22]
port 543 nsew signal output
rlabel metal2 s 42364 953270 42420 953750 6 gpio_inp_dis[23]
port 544 nsew signal output
rlabel metal3 s -424 920357 56 920427 4 gpio_inp_dis[24]
port 545 nsew signal output
rlabel metal3 s -424 750557 56 750627 4 gpio_inp_dis[25]
port 546 nsew signal output
rlabel metal3 s -424 707357 56 707427 4 gpio_inp_dis[26]
port 547 nsew signal output
rlabel metal3 s -424 664157 56 664227 4 gpio_inp_dis[27]
port 548 nsew signal output
rlabel metal3 s -424 620957 56 621027 4 gpio_inp_dis[28]
port 549 nsew signal output
rlabel metal3 s -424 577757 56 577827 4 gpio_inp_dis[29]
port 550 nsew signal output
rlabel metal3 s 633270 155699 633750 155769 6 gpio_inp_dis[2]
port 551 nsew signal output
rlabel metal3 s -424 534557 56 534627 4 gpio_inp_dis[30]
port 552 nsew signal output
rlabel metal3 s -424 491357 56 491427 4 gpio_inp_dis[31]
port 553 nsew signal output
rlabel metal3 s -424 363757 56 363827 4 gpio_inp_dis[32]
port 554 nsew signal output
rlabel metal3 s -424 320557 56 320627 4 gpio_inp_dis[33]
port 555 nsew signal output
rlabel metal3 s -424 277357 56 277427 4 gpio_inp_dis[34]
port 556 nsew signal output
rlabel metal3 s -424 234157 56 234227 4 gpio_inp_dis[35]
port 557 nsew signal output
rlabel metal3 s -424 190956 56 191028 4 gpio_inp_dis[36]
port 558 nsew signal output
rlabel metal3 s -424 147756 56 147828 4 gpio_inp_dis[37]
port 559 nsew signal output
rlabel metal2 s 151906 -424 151962 56 8 gpio_inp_dis[38]
port 560 nsew signal output
rlabel metal2 s 260506 -424 260562 56 8 gpio_inp_dis[39]
port 561 nsew signal output
rlabel metal3 s 633270 200899 633750 200969 6 gpio_inp_dis[3]
port 562 nsew signal output
rlabel metal2 s 315306 -424 315362 56 8 gpio_inp_dis[40]
port 563 nsew signal output
rlabel metal2 s 370106 -424 370162 56 8 gpio_inp_dis[41]
port 564 nsew signal output
rlabel metal2 s 424906 -424 424962 56 8 gpio_inp_dis[42]
port 565 nsew signal output
rlabel metal2 s 479706 -424 479762 56 8 gpio_inp_dis[43]
port 566 nsew signal output
rlabel metal3 s 633270 245899 633750 245969 6 gpio_inp_dis[4]
port 567 nsew signal output
rlabel metal3 s 633270 290899 633750 290969 6 gpio_inp_dis[5]
port 568 nsew signal output
rlabel metal3 s 633270 336099 633750 336169 6 gpio_inp_dis[6]
port 569 nsew signal output
rlabel metal3 s 633270 513299 633750 513369 6 gpio_inp_dis[7]
port 570 nsew signal output
rlabel metal3 s 633270 558499 633750 558569 6 gpio_inp_dis[8]
port 571 nsew signal output
rlabel metal3 s 633270 603499 633750 603569 6 gpio_inp_dis[9]
port 572 nsew signal output
rlabel metal3 s 633270 76005 633590 76067 6 gpio_loopback_one[0]
port 573 nsew signal input
rlabel metal3 s 633270 658005 633590 658067 6 gpio_loopback_one[10]
port 574 nsew signal input
rlabel metal3 s 633270 703005 633590 703067 6 gpio_loopback_one[11]
port 575 nsew signal input
rlabel metal3 s 633270 748005 633590 748067 6 gpio_loopback_one[12]
port 576 nsew signal input
rlabel metal3 s 633270 837005 633590 837067 6 gpio_loopback_one[13]
port 577 nsew signal input
rlabel metal3 s 633270 927005 633590 927067 6 gpio_loopback_one[14]
port 578 nsew signal input
rlabel metal2 s 578298 953270 578358 953590 6 gpio_loopback_one[15]
port 579 nsew signal input
rlabel metal2 s 478898 953270 478958 953590 6 gpio_loopback_one[16]
port 580 nsew signal input
rlabel metal2 s 427698 953270 427758 953590 6 gpio_loopback_one[17]
port 581 nsew signal input
rlabel metal2 s 338698 953270 338758 953590 6 gpio_loopback_one[18]
port 582 nsew signal input
rlabel metal2 s 234298 953270 234358 953590 6 gpio_loopback_one[19]
port 583 nsew signal input
rlabel metal3 s 633270 121005 633590 121067 6 gpio_loopback_one[1]
port 584 nsew signal input
rlabel metal2 s 183098 953270 183158 953590 6 gpio_loopback_one[20]
port 585 nsew signal input
rlabel metal2 s 131898 953270 131958 953590 6 gpio_loopback_one[21]
port 586 nsew signal input
rlabel metal2 s 80698 953270 80758 953590 6 gpio_loopback_one[22]
port 587 nsew signal input
rlabel metal2 s 29498 953270 29558 953590 6 gpio_loopback_one[23]
port 588 nsew signal input
rlabel metal3 s -264 906644 56 906704 4 gpio_loopback_one[24]
port 589 nsew signal input
rlabel metal3 s -264 736644 56 736704 4 gpio_loopback_one[25]
port 590 nsew signal input
rlabel metal3 s -264 693644 56 693704 4 gpio_loopback_one[26]
port 591 nsew signal input
rlabel metal3 s -264 650644 56 650704 4 gpio_loopback_one[27]
port 592 nsew signal input
rlabel metal3 s -264 607644 56 607704 4 gpio_loopback_one[28]
port 593 nsew signal input
rlabel metal3 s -264 564644 56 564704 4 gpio_loopback_one[29]
port 594 nsew signal input
rlabel metal3 s 633270 166005 633590 166067 6 gpio_loopback_one[2]
port 595 nsew signal input
rlabel metal3 s -264 521644 56 521704 4 gpio_loopback_one[30]
port 596 nsew signal input
rlabel metal3 s -264 478644 56 478704 4 gpio_loopback_one[31]
port 597 nsew signal input
rlabel metal3 s -264 349644 56 349704 4 gpio_loopback_one[32]
port 598 nsew signal input
rlabel metal3 s -264 306644 56 306704 4 gpio_loopback_one[33]
port 599 nsew signal input
rlabel metal3 s -264 263644 56 263704 4 gpio_loopback_one[34]
port 600 nsew signal input
rlabel metal3 s -264 220644 56 220704 4 gpio_loopback_one[35]
port 601 nsew signal input
rlabel metal3 s -264 177644 56 177704 4 gpio_loopback_one[36]
port 602 nsew signal input
rlabel metal3 s -264 134644 56 134704 4 gpio_loopback_one[37]
port 603 nsew signal input
rlabel metal2 s 160580 -260 160632 56 8 gpio_loopback_one[38]
port 604 nsew signal input
rlabel metal2 s 269180 -260 269232 56 8 gpio_loopback_one[39]
port 605 nsew signal input
rlabel metal3 s 633270 211005 633590 211067 6 gpio_loopback_one[3]
port 606 nsew signal input
rlabel metal2 s 323980 -260 324032 56 8 gpio_loopback_one[40]
port 607 nsew signal input
rlabel metal2 s 378780 -260 378832 56 8 gpio_loopback_one[41]
port 608 nsew signal input
rlabel metal2 s 433580 -260 433632 56 8 gpio_loopback_one[42]
port 609 nsew signal input
rlabel metal2 s 488380 -260 488432 56 8 gpio_loopback_one[43]
port 610 nsew signal input
rlabel metal3 s 633270 256005 633590 256067 6 gpio_loopback_one[4]
port 611 nsew signal input
rlabel metal3 s 633270 301005 633590 301067 6 gpio_loopback_one[5]
port 612 nsew signal input
rlabel metal3 s 633270 346005 633590 346067 6 gpio_loopback_one[6]
port 613 nsew signal input
rlabel metal3 s 633270 523005 633590 523067 6 gpio_loopback_one[7]
port 614 nsew signal input
rlabel metal3 s 633270 568005 633590 568067 6 gpio_loopback_one[8]
port 615 nsew signal input
rlabel metal3 s 633270 613005 633590 613067 6 gpio_loopback_one[9]
port 616 nsew signal input
rlabel metal3 s 633270 78007 633590 78069 6 gpio_loopback_zero[0]
port 617 nsew signal input
rlabel metal3 s 633270 660007 633590 660069 6 gpio_loopback_zero[10]
port 618 nsew signal input
rlabel metal3 s 633270 705007 633590 705069 6 gpio_loopback_zero[11]
port 619 nsew signal input
rlabel metal3 s 633270 750007 633590 750069 6 gpio_loopback_zero[12]
port 620 nsew signal input
rlabel metal3 s 633270 839007 633590 839069 6 gpio_loopback_zero[13]
port 621 nsew signal input
rlabel metal3 s 633270 929007 633590 929069 6 gpio_loopback_zero[14]
port 622 nsew signal input
rlabel metal2 s 576298 953270 576358 953590 6 gpio_loopback_zero[15]
port 623 nsew signal input
rlabel metal2 s 476898 953270 476958 953590 6 gpio_loopback_zero[16]
port 624 nsew signal input
rlabel metal2 s 425698 953270 425758 953590 6 gpio_loopback_zero[17]
port 625 nsew signal input
rlabel metal2 s 336698 953270 336758 953590 6 gpio_loopback_zero[18]
port 626 nsew signal input
rlabel metal2 s 232298 953270 232358 953590 6 gpio_loopback_zero[19]
port 627 nsew signal input
rlabel metal3 s 633270 123007 633590 123069 6 gpio_loopback_zero[1]
port 628 nsew signal input
rlabel metal2 s 181098 953270 181158 953590 6 gpio_loopback_zero[20]
port 629 nsew signal input
rlabel metal2 s 129898 953270 129958 953590 6 gpio_loopback_zero[21]
port 630 nsew signal input
rlabel metal2 s 78698 953270 78758 953590 6 gpio_loopback_zero[22]
port 631 nsew signal input
rlabel metal2 s 27498 953270 27558 953590 6 gpio_loopback_zero[23]
port 632 nsew signal input
rlabel metal3 s -264 904644 56 904704 4 gpio_loopback_zero[24]
port 633 nsew signal input
rlabel metal3 s -264 734644 56 734704 4 gpio_loopback_zero[25]
port 634 nsew signal input
rlabel metal3 s -264 691644 56 691704 4 gpio_loopback_zero[26]
port 635 nsew signal input
rlabel metal3 s -264 648644 56 648704 4 gpio_loopback_zero[27]
port 636 nsew signal input
rlabel metal3 s -264 605644 56 605704 4 gpio_loopback_zero[28]
port 637 nsew signal input
rlabel metal3 s -264 562644 56 562704 4 gpio_loopback_zero[29]
port 638 nsew signal input
rlabel metal3 s 633270 168007 633590 168069 6 gpio_loopback_zero[2]
port 639 nsew signal input
rlabel metal3 s -264 519644 56 519704 4 gpio_loopback_zero[30]
port 640 nsew signal input
rlabel metal3 s -264 476644 56 476704 4 gpio_loopback_zero[31]
port 641 nsew signal input
rlabel metal3 s -264 347644 56 347704 4 gpio_loopback_zero[32]
port 642 nsew signal input
rlabel metal3 s -264 304644 56 304704 4 gpio_loopback_zero[33]
port 643 nsew signal input
rlabel metal3 s -264 261644 56 261704 4 gpio_loopback_zero[34]
port 644 nsew signal input
rlabel metal3 s -264 218644 56 218704 4 gpio_loopback_zero[35]
port 645 nsew signal input
rlabel metal3 s -264 175644 56 175704 4 gpio_loopback_zero[36]
port 646 nsew signal input
rlabel metal3 s -264 132644 56 132704 4 gpio_loopback_zero[37]
port 647 nsew signal input
rlabel metal2 s 163791 -259 163843 57 8 gpio_loopback_zero[38]
port 648 nsew signal input
rlabel metal2 s 273360 -260 273412 56 8 gpio_loopback_zero[39]
port 649 nsew signal input
rlabel metal3 s 633270 213007 633590 213069 6 gpio_loopback_zero[3]
port 650 nsew signal input
rlabel metal2 s 328165 -282 328217 34 8 gpio_loopback_zero[40]
port 651 nsew signal input
rlabel metal2 s 382978 -260 383030 56 8 gpio_loopback_zero[41]
port 652 nsew signal input
rlabel metal2 s 437778 -260 437830 56 8 gpio_loopback_zero[42]
port 653 nsew signal input
rlabel metal2 s 492635 -260 492687 56 8 gpio_loopback_zero[43]
port 654 nsew signal input
rlabel metal3 s 633270 258007 633590 258069 6 gpio_loopback_zero[4]
port 655 nsew signal input
rlabel metal3 s 633270 303007 633590 303069 6 gpio_loopback_zero[5]
port 656 nsew signal input
rlabel metal3 s 633270 348007 633590 348069 6 gpio_loopback_zero[6]
port 657 nsew signal input
rlabel metal3 s 633270 525007 633590 525069 6 gpio_loopback_zero[7]
port 658 nsew signal input
rlabel metal3 s 633270 570007 633590 570069 6 gpio_loopback_zero[8]
port 659 nsew signal input
rlabel metal3 s 633270 615007 633590 615069 6 gpio_loopback_zero[9]
port 660 nsew signal input
rlabel metal3 s 633270 72951 633750 73021 6 gpio_oeb[0]
port 661 nsew signal output
rlabel metal3 s 633270 656151 633750 656221 6 gpio_oeb[10]
port 662 nsew signal output
rlabel metal3 s 633270 701151 633750 701221 6 gpio_oeb[11]
port 663 nsew signal output
rlabel metal3 s 633270 746151 633750 746221 6 gpio_oeb[12]
port 664 nsew signal output
rlabel metal3 s 633270 835351 633750 835421 6 gpio_oeb[13]
port 665 nsew signal output
rlabel metal3 s 633270 924551 633750 924621 6 gpio_oeb[14]
port 666 nsew signal output
rlabel metal2 s 584712 953270 584768 953750 6 gpio_oeb[15]
port 667 nsew signal output
rlabel metal2 s 482912 953270 482968 953750 6 gpio_oeb[16]
port 668 nsew signal output
rlabel metal2 s 431512 953270 431568 953750 6 gpio_oeb[17]
port 669 nsew signal output
rlabel metal2 s 342512 953270 342568 953750 6 gpio_oeb[18]
port 670 nsew signal output
rlabel metal2 s 240712 953270 240768 953750 6 gpio_oeb[19]
port 671 nsew signal output
rlabel metal3 s 633270 118151 633750 118221 6 gpio_oeb[1]
port 672 nsew signal output
rlabel metal2 s 189112 953270 189168 953750 6 gpio_oeb[20]
port 673 nsew signal output
rlabel metal2 s 137712 953270 137768 953750 6 gpio_oeb[21]
port 674 nsew signal output
rlabel metal2 s 86312 953270 86368 953750 6 gpio_oeb[22]
port 675 nsew signal output
rlabel metal2 s 34912 953270 34968 953750 6 gpio_oeb[23]
port 676 nsew signal output
rlabel metal3 s -424 912905 56 912975 4 gpio_oeb[24]
port 677 nsew signal output
rlabel metal3 s -424 743105 56 743175 4 gpio_oeb[25]
port 678 nsew signal output
rlabel metal3 s -424 699905 56 699975 4 gpio_oeb[26]
port 679 nsew signal output
rlabel metal3 s -424 656705 56 656775 4 gpio_oeb[27]
port 680 nsew signal output
rlabel metal3 s -424 613505 56 613575 4 gpio_oeb[28]
port 681 nsew signal output
rlabel metal3 s -424 570305 56 570375 4 gpio_oeb[29]
port 682 nsew signal output
rlabel metal3 s 633270 163151 633750 163221 6 gpio_oeb[2]
port 683 nsew signal output
rlabel metal3 s -424 527105 56 527175 4 gpio_oeb[30]
port 684 nsew signal output
rlabel metal3 s -424 483905 56 483975 4 gpio_oeb[31]
port 685 nsew signal output
rlabel metal3 s -424 356305 56 356375 4 gpio_oeb[32]
port 686 nsew signal output
rlabel metal3 s -424 313105 56 313175 4 gpio_oeb[33]
port 687 nsew signal output
rlabel metal3 s -424 269905 56 269975 4 gpio_oeb[34]
port 688 nsew signal output
rlabel metal3 s -424 226705 56 226775 4 gpio_oeb[35]
port 689 nsew signal output
rlabel metal3 s -424 183504 56 183576 4 gpio_oeb[36]
port 690 nsew signal output
rlabel metal3 s -424 140304 56 140376 4 gpio_oeb[37]
port 691 nsew signal output
rlabel metal2 s 159358 -424 159414 56 8 gpio_oeb[38]
port 692 nsew signal output
rlabel metal2 s 267958 -424 268014 56 8 gpio_oeb[39]
port 693 nsew signal output
rlabel metal3 s 633270 208351 633750 208421 6 gpio_oeb[3]
port 694 nsew signal output
rlabel metal2 s 322758 -424 322814 56 8 gpio_oeb[40]
port 695 nsew signal output
rlabel metal2 s 377558 -424 377614 56 8 gpio_oeb[41]
port 696 nsew signal output
rlabel metal2 s 432358 -424 432414 56 8 gpio_oeb[42]
port 697 nsew signal output
rlabel metal2 s 487158 -424 487214 56 8 gpio_oeb[43]
port 698 nsew signal output
rlabel metal3 s 633270 253351 633750 253421 6 gpio_oeb[4]
port 699 nsew signal output
rlabel metal3 s 633270 298351 633750 298421 6 gpio_oeb[5]
port 700 nsew signal output
rlabel metal3 s 633270 343551 633750 343621 6 gpio_oeb[6]
port 701 nsew signal output
rlabel metal3 s 633270 520751 633750 520821 6 gpio_oeb[7]
port 702 nsew signal output
rlabel metal3 s 633270 565951 633750 566021 6 gpio_oeb[8]
port 703 nsew signal output
rlabel metal3 s 633270 610951 633750 611021 6 gpio_oeb[9]
port 704 nsew signal output
rlabel metal3 s 633270 69823 633750 69893 6 gpio_out[0]
port 705 nsew signal output
rlabel metal3 s 633270 653023 633750 653093 6 gpio_out[10]
port 706 nsew signal output
rlabel metal3 s 633270 698023 633750 698093 6 gpio_out[11]
port 707 nsew signal output
rlabel metal3 s 633270 743023 633750 743093 6 gpio_out[12]
port 708 nsew signal output
rlabel metal3 s 633270 832223 633750 832293 6 gpio_out[13]
port 709 nsew signal output
rlabel metal3 s 633270 921423 633750 921493 6 gpio_out[14]
port 710 nsew signal output
rlabel metal2 s 587840 953270 587896 953750 6 gpio_out[15]
port 711 nsew signal output
rlabel metal2 s 486040 953270 486096 953750 6 gpio_out[16]
port 712 nsew signal output
rlabel metal2 s 434640 953270 434696 953750 6 gpio_out[17]
port 713 nsew signal output
rlabel metal2 s 345640 953270 345696 953750 6 gpio_out[18]
port 714 nsew signal output
rlabel metal2 s 243840 953270 243896 953750 6 gpio_out[19]
port 715 nsew signal output
rlabel metal3 s 633270 115023 633750 115093 6 gpio_out[1]
port 716 nsew signal output
rlabel metal2 s 192240 953270 192296 953750 6 gpio_out[20]
port 717 nsew signal output
rlabel metal2 s 140840 953270 140896 953750 6 gpio_out[21]
port 718 nsew signal output
rlabel metal2 s 89440 953270 89496 953750 6 gpio_out[22]
port 719 nsew signal output
rlabel metal2 s 38040 953270 38096 953750 6 gpio_out[23]
port 720 nsew signal output
rlabel metal3 s -424 916033 56 916103 4 gpio_out[24]
port 721 nsew signal output
rlabel metal3 s -424 746233 56 746303 4 gpio_out[25]
port 722 nsew signal output
rlabel metal3 s -424 703033 56 703103 4 gpio_out[26]
port 723 nsew signal output
rlabel metal3 s -424 659833 56 659903 4 gpio_out[27]
port 724 nsew signal output
rlabel metal3 s -424 616633 56 616703 4 gpio_out[28]
port 725 nsew signal output
rlabel metal3 s -424 573433 56 573503 4 gpio_out[29]
port 726 nsew signal output
rlabel metal3 s 633270 160023 633750 160093 6 gpio_out[2]
port 727 nsew signal output
rlabel metal3 s -424 530233 56 530303 4 gpio_out[30]
port 728 nsew signal output
rlabel metal3 s -424 487033 56 487103 4 gpio_out[31]
port 729 nsew signal output
rlabel metal3 s -424 359433 56 359503 4 gpio_out[32]
port 730 nsew signal output
rlabel metal3 s -424 316233 56 316303 4 gpio_out[33]
port 731 nsew signal output
rlabel metal3 s -424 273033 56 273103 4 gpio_out[34]
port 732 nsew signal output
rlabel metal3 s -424 229833 56 229903 4 gpio_out[35]
port 733 nsew signal output
rlabel metal3 s -424 186632 56 186704 4 gpio_out[36]
port 734 nsew signal output
rlabel metal3 s -424 143432 56 143504 4 gpio_out[37]
port 735 nsew signal output
rlabel metal2 s 156230 -424 156286 56 8 gpio_out[38]
port 736 nsew signal output
rlabel metal2 s 264830 -424 264886 56 8 gpio_out[39]
port 737 nsew signal output
rlabel metal3 s 633270 205223 633750 205293 6 gpio_out[3]
port 738 nsew signal output
rlabel metal2 s 319630 -424 319686 56 8 gpio_out[40]
port 739 nsew signal output
rlabel metal2 s 374430 -424 374486 56 8 gpio_out[41]
port 740 nsew signal output
rlabel metal2 s 429230 -424 429286 56 8 gpio_out[42]
port 741 nsew signal output
rlabel metal2 s 484030 -424 484086 56 8 gpio_out[43]
port 742 nsew signal output
rlabel metal3 s 633270 250223 633750 250293 6 gpio_out[4]
port 743 nsew signal output
rlabel metal3 s 633270 295223 633750 295293 6 gpio_out[5]
port 744 nsew signal output
rlabel metal3 s 633270 340423 633750 340493 6 gpio_out[6]
port 745 nsew signal output
rlabel metal3 s 633270 517623 633750 517693 6 gpio_out[7]
port 746 nsew signal output
rlabel metal3 s 633270 562823 633750 562893 6 gpio_out[8]
port 747 nsew signal output
rlabel metal3 s 633270 607823 633750 607893 6 gpio_out[9]
port 748 nsew signal output
rlabel metal3 s 633270 60623 633750 60693 6 gpio_slow_sel[0]
port 749 nsew signal output
rlabel metal3 s 633270 643823 633750 643893 6 gpio_slow_sel[10]
port 750 nsew signal output
rlabel metal3 s 633270 688823 633750 688893 6 gpio_slow_sel[11]
port 751 nsew signal output
rlabel metal3 s 633270 733823 633750 733893 6 gpio_slow_sel[12]
port 752 nsew signal output
rlabel metal3 s 633270 823023 633750 823093 6 gpio_slow_sel[13]
port 753 nsew signal output
rlabel metal3 s 633270 912223 633750 912293 6 gpio_slow_sel[14]
port 754 nsew signal output
rlabel metal2 s 597040 953270 597096 953750 6 gpio_slow_sel[15]
port 755 nsew signal output
rlabel metal2 s 495240 953270 495296 953750 6 gpio_slow_sel[16]
port 756 nsew signal output
rlabel metal2 s 443840 953270 443896 953750 6 gpio_slow_sel[17]
port 757 nsew signal output
rlabel metal2 s 354840 953270 354896 953750 6 gpio_slow_sel[18]
port 758 nsew signal output
rlabel metal2 s 253040 953270 253096 953750 6 gpio_slow_sel[19]
port 759 nsew signal output
rlabel metal3 s 633270 105823 633750 105893 6 gpio_slow_sel[1]
port 760 nsew signal output
rlabel metal2 s 201440 953270 201496 953750 6 gpio_slow_sel[20]
port 761 nsew signal output
rlabel metal2 s 150040 953270 150096 953750 6 gpio_slow_sel[21]
port 762 nsew signal output
rlabel metal2 s 98640 953270 98696 953750 6 gpio_slow_sel[22]
port 763 nsew signal output
rlabel metal2 s 47240 953270 47296 953750 6 gpio_slow_sel[23]
port 764 nsew signal output
rlabel metal3 s -424 925233 56 925303 4 gpio_slow_sel[24]
port 765 nsew signal output
rlabel metal3 s -424 755433 56 755503 4 gpio_slow_sel[25]
port 766 nsew signal output
rlabel metal3 s -424 712233 56 712303 4 gpio_slow_sel[26]
port 767 nsew signal output
rlabel metal3 s -424 669033 56 669103 4 gpio_slow_sel[27]
port 768 nsew signal output
rlabel metal3 s -424 625833 56 625903 4 gpio_slow_sel[28]
port 769 nsew signal output
rlabel metal3 s -424 582633 56 582703 4 gpio_slow_sel[29]
port 770 nsew signal output
rlabel metal3 s 633270 150823 633750 150893 6 gpio_slow_sel[2]
port 771 nsew signal output
rlabel metal3 s -424 539433 56 539503 4 gpio_slow_sel[30]
port 772 nsew signal output
rlabel metal3 s -424 496233 56 496303 4 gpio_slow_sel[31]
port 773 nsew signal output
rlabel metal3 s -424 368633 56 368703 4 gpio_slow_sel[32]
port 774 nsew signal output
rlabel metal3 s -424 325433 56 325503 4 gpio_slow_sel[33]
port 775 nsew signal output
rlabel metal3 s -424 282233 56 282303 4 gpio_slow_sel[34]
port 776 nsew signal output
rlabel metal3 s -424 239033 56 239103 4 gpio_slow_sel[35]
port 777 nsew signal output
rlabel metal3 s -424 195832 56 195904 4 gpio_slow_sel[36]
port 778 nsew signal output
rlabel metal3 s -424 152632 56 152704 4 gpio_slow_sel[37]
port 779 nsew signal output
rlabel metal2 s 147030 -424 147086 56 8 gpio_slow_sel[38]
port 780 nsew signal output
rlabel metal2 s 255630 -424 255686 56 8 gpio_slow_sel[39]
port 781 nsew signal output
rlabel metal3 s 633270 196023 633750 196093 6 gpio_slow_sel[3]
port 782 nsew signal output
rlabel metal2 s 310430 -424 310486 56 8 gpio_slow_sel[40]
port 783 nsew signal output
rlabel metal2 s 365230 -424 365286 56 8 gpio_slow_sel[41]
port 784 nsew signal output
rlabel metal2 s 420030 -424 420086 56 8 gpio_slow_sel[42]
port 785 nsew signal output
rlabel metal2 s 474830 -424 474886 56 8 gpio_slow_sel[43]
port 786 nsew signal output
rlabel metal3 s 633270 241023 633750 241093 6 gpio_slow_sel[4]
port 787 nsew signal output
rlabel metal3 s 633270 286023 633750 286093 6 gpio_slow_sel[5]
port 788 nsew signal output
rlabel metal3 s 633270 331223 633750 331293 6 gpio_slow_sel[6]
port 789 nsew signal output
rlabel metal3 s 633270 508423 633750 508493 6 gpio_slow_sel[7]
port 790 nsew signal output
rlabel metal3 s 633270 553623 633750 553693 6 gpio_slow_sel[8]
port 791 nsew signal output
rlabel metal3 s 633270 598623 633750 598693 6 gpio_slow_sel[9]
port 792 nsew signal output
rlabel metal3 s 633270 71663 633750 71733 6 gpio_vtrip_sel[0]
port 793 nsew signal output
rlabel metal3 s 633270 654863 633750 654933 6 gpio_vtrip_sel[10]
port 794 nsew signal output
rlabel metal3 s 633270 699863 633750 699933 6 gpio_vtrip_sel[11]
port 795 nsew signal output
rlabel metal3 s 633270 744863 633750 744933 6 gpio_vtrip_sel[12]
port 796 nsew signal output
rlabel metal3 s 633270 834063 633750 834133 6 gpio_vtrip_sel[13]
port 797 nsew signal output
rlabel metal3 s 633270 923263 633750 923333 6 gpio_vtrip_sel[14]
port 798 nsew signal output
rlabel metal2 s 586000 953270 586056 953750 6 gpio_vtrip_sel[15]
port 799 nsew signal output
rlabel metal2 s 484200 953270 484256 953750 6 gpio_vtrip_sel[16]
port 800 nsew signal output
rlabel metal2 s 432800 953270 432856 953750 6 gpio_vtrip_sel[17]
port 801 nsew signal output
rlabel metal2 s 343800 953270 343856 953750 6 gpio_vtrip_sel[18]
port 802 nsew signal output
rlabel metal2 s 242000 953270 242056 953750 6 gpio_vtrip_sel[19]
port 803 nsew signal output
rlabel metal3 s 633270 116863 633750 116933 6 gpio_vtrip_sel[1]
port 804 nsew signal output
rlabel metal2 s 190400 953270 190456 953750 6 gpio_vtrip_sel[20]
port 805 nsew signal output
rlabel metal2 s 139000 953270 139056 953750 6 gpio_vtrip_sel[21]
port 806 nsew signal output
rlabel metal2 s 87600 953270 87656 953750 6 gpio_vtrip_sel[22]
port 807 nsew signal output
rlabel metal2 s 36200 953270 36256 953750 6 gpio_vtrip_sel[23]
port 808 nsew signal output
rlabel metal3 s -424 914193 56 914263 4 gpio_vtrip_sel[24]
port 809 nsew signal output
rlabel metal3 s -424 744393 56 744463 4 gpio_vtrip_sel[25]
port 810 nsew signal output
rlabel metal3 s -424 701193 56 701263 4 gpio_vtrip_sel[26]
port 811 nsew signal output
rlabel metal3 s -424 657993 56 658063 4 gpio_vtrip_sel[27]
port 812 nsew signal output
rlabel metal3 s -424 614793 56 614863 4 gpio_vtrip_sel[28]
port 813 nsew signal output
rlabel metal3 s -424 571593 56 571663 4 gpio_vtrip_sel[29]
port 814 nsew signal output
rlabel metal3 s 633270 161863 633750 161933 6 gpio_vtrip_sel[2]
port 815 nsew signal output
rlabel metal3 s -424 528393 56 528463 4 gpio_vtrip_sel[30]
port 816 nsew signal output
rlabel metal3 s -424 485193 56 485263 4 gpio_vtrip_sel[31]
port 817 nsew signal output
rlabel metal3 s -424 357593 56 357663 4 gpio_vtrip_sel[32]
port 818 nsew signal output
rlabel metal3 s -424 314393 56 314463 4 gpio_vtrip_sel[33]
port 819 nsew signal output
rlabel metal3 s -424 271193 56 271263 4 gpio_vtrip_sel[34]
port 820 nsew signal output
rlabel metal3 s -424 227993 56 228063 4 gpio_vtrip_sel[35]
port 821 nsew signal output
rlabel metal3 s -424 184792 56 184864 4 gpio_vtrip_sel[36]
port 822 nsew signal output
rlabel metal3 s -424 141592 56 141664 4 gpio_vtrip_sel[37]
port 823 nsew signal output
rlabel metal2 s 158070 -424 158126 56 8 gpio_vtrip_sel[38]
port 824 nsew signal output
rlabel metal2 s 266670 -424 266726 56 8 gpio_vtrip_sel[39]
port 825 nsew signal output
rlabel metal3 s 633270 207063 633750 207133 6 gpio_vtrip_sel[3]
port 826 nsew signal output
rlabel metal2 s 321470 -424 321526 56 8 gpio_vtrip_sel[40]
port 827 nsew signal output
rlabel metal2 s 376270 -424 376326 56 8 gpio_vtrip_sel[41]
port 828 nsew signal output
rlabel metal2 s 431070 -424 431126 56 8 gpio_vtrip_sel[42]
port 829 nsew signal output
rlabel metal2 s 485870 -424 485926 56 8 gpio_vtrip_sel[43]
port 830 nsew signal output
rlabel metal3 s 633270 252063 633750 252133 6 gpio_vtrip_sel[4]
port 831 nsew signal output
rlabel metal3 s 633270 297063 633750 297133 6 gpio_vtrip_sel[5]
port 832 nsew signal output
rlabel metal3 s 633270 342263 633750 342333 6 gpio_vtrip_sel[6]
port 833 nsew signal output
rlabel metal3 s 633270 519463 633750 519533 6 gpio_vtrip_sel[7]
port 834 nsew signal output
rlabel metal3 s 633270 564663 633750 564733 6 gpio_vtrip_sel[8]
port 835 nsew signal output
rlabel metal3 s 633270 609663 633750 609733 6 gpio_vtrip_sel[9]
port 836 nsew signal output
rlabel metal2 s 605082 -260 605134 56 8 mask_rev[0]
port 837 nsew signal input
rlabel metal2 s 607322 -260 607374 56 8 mask_rev[10]
port 838 nsew signal input
rlabel metal2 s 607546 -260 607598 56 8 mask_rev[11]
port 839 nsew signal input
rlabel metal2 s 607770 -260 607822 56 8 mask_rev[12]
port 840 nsew signal input
rlabel metal2 s 607994 -260 608046 56 8 mask_rev[13]
port 841 nsew signal input
rlabel metal2 s 608218 -260 608270 56 8 mask_rev[14]
port 842 nsew signal input
rlabel metal2 s 608442 -260 608494 56 8 mask_rev[15]
port 843 nsew signal input
rlabel metal2 s 608666 -260 608718 56 8 mask_rev[16]
port 844 nsew signal input
rlabel metal2 s 608890 -260 608942 56 8 mask_rev[17]
port 845 nsew signal input
rlabel metal2 s 609114 -260 609166 56 8 mask_rev[18]
port 846 nsew signal input
rlabel metal2 s 609338 -260 609390 56 8 mask_rev[19]
port 847 nsew signal input
rlabel metal2 s 605306 -260 605358 56 8 mask_rev[1]
port 848 nsew signal input
rlabel metal2 s 609562 -260 609614 56 8 mask_rev[20]
port 849 nsew signal input
rlabel metal2 s 609786 -260 609838 56 8 mask_rev[21]
port 850 nsew signal input
rlabel metal2 s 610010 -260 610062 56 8 mask_rev[22]
port 851 nsew signal input
rlabel metal2 s 610234 -260 610286 56 8 mask_rev[23]
port 852 nsew signal input
rlabel metal2 s 610458 -260 610510 56 8 mask_rev[24]
port 853 nsew signal input
rlabel metal2 s 610682 -260 610734 56 8 mask_rev[25]
port 854 nsew signal input
rlabel metal2 s 610906 -260 610958 56 8 mask_rev[26]
port 855 nsew signal input
rlabel metal2 s 611130 -260 611182 56 8 mask_rev[27]
port 856 nsew signal input
rlabel metal2 s 611354 -260 611406 56 8 mask_rev[28]
port 857 nsew signal input
rlabel metal2 s 611578 -260 611630 56 8 mask_rev[29]
port 858 nsew signal input
rlabel metal2 s 605530 -260 605582 56 8 mask_rev[2]
port 859 nsew signal input
rlabel metal2 s 611802 -260 611854 56 8 mask_rev[30]
port 860 nsew signal input
rlabel metal2 s 612026 -260 612078 56 8 mask_rev[31]
port 861 nsew signal input
rlabel metal2 s 605754 -260 605806 56 8 mask_rev[3]
port 862 nsew signal input
rlabel metal2 s 605978 -260 606030 56 8 mask_rev[4]
port 863 nsew signal input
rlabel metal2 s 606202 -260 606254 56 8 mask_rev[5]
port 864 nsew signal input
rlabel metal2 s 606426 -260 606478 56 8 mask_rev[6]
port 865 nsew signal input
rlabel metal2 s 606650 -260 606702 56 8 mask_rev[7]
port 866 nsew signal input
rlabel metal2 s 606874 -260 606926 56 8 mask_rev[8]
port 867 nsew signal input
rlabel metal2 s 607098 -260 607150 56 8 mask_rev[9]
port 868 nsew signal input
rlabel metal3 s -284 53372 56 53442 4 por_l
port 869 nsew signal input
rlabel metal3 s -284 53147 56 53217 4 porb_h
port 870 nsew signal input
rlabel metal3 s -284 53595 56 53665 4 porb_l
port 871 nsew signal input
rlabel metal2 s 99571 -90 99637 56 8 resetb_h
port 872 nsew signal input
rlabel metal2 s 110164 -116 110220 56 8 resetb_l
port 873 nsew signal input
rlabel metal4 s 4804 4960 8804 948128 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 4804 4960 628524 8960 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 4804 944128 628524 948128 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 624524 4960 628524 948128 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 11050 480 12330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 19050 480 20330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 27050 480 28330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 35050 480 36330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 43050 480 44330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 51050 480 52330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 59050 480 60330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 67050 480 68330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 75050 480 76330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 83050 480 84330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 91050 480 92330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 91050 709904 92330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 99050 480 100330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 99050 709904 100330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 107050 480 108330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 107050 709904 108330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 115050 480 116330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 115050 709904 116330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 123050 480 124330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 123050 709904 124330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 131050 480 132330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 131050 709904 132330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 139050 480 140330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 139050 709904 140330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 147050 480 148330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 147050 709904 148330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 155050 480 156330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 155050 709904 156330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 163050 480 164330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 163050 709904 164330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 171050 480 172330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 171050 709904 172330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 179050 480 180330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 179050 709904 180330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 187050 480 188330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 187050 709904 188330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 195050 480 196330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 195050 709904 196330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 203050 480 204330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 203050 709904 204330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 211050 480 212330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 211050 709904 212330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 219050 480 220330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 219050 709904 220330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 227050 480 228330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 227050 709904 228330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 235050 480 236330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 235050 709904 236330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 243050 480 244330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 243050 709904 244330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 251050 480 252330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 251050 709904 252330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 259050 480 260330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 259050 709904 260330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 267050 480 268330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 267050 709904 268330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 275050 480 276330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 275050 709904 276330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 283050 480 284330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 283050 709904 284330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 291050 480 292330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 291050 709904 292330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 299050 480 300330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 299050 709904 300330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 307050 480 308330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 307050 709904 308330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 315050 480 316330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 315050 709904 316330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 323050 480 324330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 323050 709904 324330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 331050 480 332330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 331050 709904 332330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 339050 480 340330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 339050 709904 340330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 347050 480 348330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 347050 709904 348330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 355050 480 356330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 355050 709904 356330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 363050 480 364330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 363050 709904 364330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 371050 480 372330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 371050 709904 372330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 379050 480 380330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 379050 709904 380330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 387050 480 388330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 387050 709904 388330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 395050 480 396330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 395050 709904 396330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 403050 480 404330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 403050 709904 404330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 411050 480 412330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 411050 709904 412330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 419050 480 420330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 419050 709904 420330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 427050 480 428330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 427050 709904 428330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 435050 480 436330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 435050 709904 436330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 443050 480 444330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 443050 709904 444330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 451050 480 452330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 451050 709904 452330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 459050 480 460330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 459050 709904 460330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 467050 480 468330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 467050 709904 468330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 475050 480 476330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 475050 709904 476330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 483050 480 484330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 483050 709904 484330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 491050 480 492330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 491050 709904 492330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 499050 480 500330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 499050 709904 500330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 507050 480 508330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 507050 709904 508330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 515050 480 516330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 515050 709904 516330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 523050 480 524330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 523050 709904 524330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 531050 480 532330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 531050 709904 532330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 539050 480 540330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 539050 709904 540330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 547050 480 548330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 547050 709904 548330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 555050 480 556330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 555050 709904 556330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 563050 480 564330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 563050 709904 564330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 571050 480 572330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 571050 709904 572330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 579050 480 580330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 579050 709904 580330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 587050 480 588330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 587050 709904 588330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 595050 480 596330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 595050 709904 596330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 603050 480 604330 389968 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 603050 709904 604330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 611050 480 612330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 619050 480 620330 952608 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 12086 633004 13366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 20086 633004 21366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 28086 633004 29366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 36086 633004 37366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 44086 633004 45366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 52086 633004 53366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 60086 633004 61366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 68086 633004 69366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 76086 633004 77366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 84086 633004 85366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 92086 633004 93366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 100086 633004 101366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 108086 633004 109366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 116086 633004 117366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 124086 633004 125366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 132086 633004 133366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 140086 633004 141366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 148086 633004 149366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 156086 633004 157366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 164086 633004 165366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 172086 633004 173366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 180086 633004 181366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 188086 633004 189366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 196086 633004 197366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 204086 633004 205366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 212086 633004 213366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 220086 633004 221366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 228086 633004 229366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 236086 633004 237366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 244086 633004 245366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 252086 633004 253366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 260086 633004 261366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 268086 633004 269366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 276086 633004 277366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 284086 633004 285366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 292086 633004 293366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 300086 633004 301366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 308086 633004 309366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 316086 633004 317366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 324086 633004 325366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 332086 633004 333366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 340086 633004 341366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 348086 633004 349366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 356086 633004 357366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 364086 633004 365366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 372086 633004 373366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 380086 633004 381366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 388086 633004 389366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 396086 633004 397366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 404086 633004 405366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 412086 633004 413366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 420086 633004 421366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 428086 633004 429366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 436086 633004 437366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 444086 633004 445366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 452086 139548 453366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 460086 139548 461366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 468086 139548 469366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 476086 139548 477366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 484086 139548 485366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 492086 139548 493366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 500086 139548 501366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 508086 139548 509366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 516086 139548 517366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 524086 139548 525366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 532086 139548 533366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 540086 139548 541366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 548086 633004 549366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 556086 633004 557366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 564086 633004 565366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 572086 633004 573366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 580086 633004 581366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 588086 633004 589366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 596086 633004 597366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 604086 633004 605366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 612086 633004 613366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 620086 633004 621366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 628086 633004 629366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 636086 633004 637366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 644086 633004 645366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 652086 633004 653366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 660086 633004 661366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 668086 633004 669366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 676086 633004 677366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 684086 633004 685366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 692086 633004 693366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 700086 633004 701366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 708086 633004 709366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 716086 633004 717366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 724086 633004 725366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 732086 633004 733366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 740086 633004 741366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 748086 633004 749366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 756086 633004 757366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 764086 633004 765366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 772086 633004 773366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 780086 633004 781366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 788086 633004 789366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 796086 633004 797366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 804086 633004 805366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 812086 633004 813366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 820086 633004 821366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 828086 633004 829366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 836086 633004 837366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 844086 633004 845366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 852086 633004 853366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 860086 633004 861366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 868086 633004 869366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 876086 633004 877366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 884086 633004 885366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 892086 633004 893366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 900086 633004 901366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 908086 633004 909366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 916086 633004 917366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 924086 633004 925366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 932086 633004 933366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 324 940086 633004 941366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 452086 633004 453366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 460086 633004 461366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 468086 633004 469366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 476086 633004 477366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 484086 633004 485366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 492086 633004 493366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 500086 633004 501366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 508086 633004 509366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 516086 633004 517366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 524086 633004 525366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 532086 633004 533366 6 vccd1
port 874 nsew power bidirectional
rlabel metal5 s 433660 540086 633004 541366 6 vccd1
port 874 nsew power bidirectional
rlabel metal4 s 324 480 4324 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 480 633004 4480 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 948608 633004 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 629004 480 633004 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 12970 480 14250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 20970 480 22250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 28970 480 30250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 36970 480 38250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 44970 480 46250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 52970 480 54250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 60970 480 62250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 68970 480 70250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 76970 480 78250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 84970 480 86250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 92970 480 94250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 92970 709904 94250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 100970 480 102250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 100970 709904 102250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 108970 480 110250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 108970 709904 110250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 116970 480 118250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 116970 709904 118250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 124970 480 126250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 124970 709904 126250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 132970 480 134250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 132970 709904 134250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 140970 480 142250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 140970 709904 142250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 148970 480 150250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 148970 709904 150250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 156970 480 158250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 156970 709904 158250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 164970 480 166250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 164970 709904 166250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 172970 480 174250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 172970 709904 174250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 180970 480 182250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 180970 709904 182250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 188970 480 190250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 188970 709904 190250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 196970 480 198250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 196970 709904 198250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 204970 480 206250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 204970 709904 206250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 212970 480 214250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 212970 709904 214250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 220970 480 222250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 220970 709904 222250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 228970 480 230250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 228970 709904 230250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 236970 480 238250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 236970 709904 238250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 244970 480 246250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 244970 709904 246250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 252970 480 254250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 252970 709904 254250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 260970 480 262250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 260970 709904 262250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 268970 480 270250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 268970 709904 270250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 276970 480 278250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 276970 709904 278250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 284970 480 286250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 284970 709904 286250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 292970 480 294250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 292970 709904 294250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 300970 480 302250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 300970 709904 302250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 308970 480 310250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 308970 709904 310250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 316970 480 318250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 316970 709904 318250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 324970 480 326250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 324970 709904 326250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 332970 480 334250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 332970 709904 334250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 340970 480 342250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 340970 709904 342250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 348970 480 350250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 348970 709904 350250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 356970 480 358250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 356970 709904 358250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 364970 480 366250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 364970 709904 366250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 372970 480 374250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 372970 709904 374250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 380970 480 382250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 380970 709904 382250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 388970 480 390250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 388970 709904 390250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 396970 480 398250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 396970 709904 398250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 404970 480 406250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 404970 709904 406250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 412970 480 414250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 412970 709904 414250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 420970 480 422250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 420970 709904 422250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 428970 480 430250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 428970 709904 430250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 436970 480 438250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 436970 709904 438250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 444970 480 446250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 444970 709904 446250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 452970 480 454250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 452970 709904 454250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 460970 480 462250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 460970 709904 462250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 468970 480 470250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 468970 709904 470250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 476970 480 478250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 476970 709904 478250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 484970 480 486250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 484970 709904 486250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 492970 480 494250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 492970 709904 494250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 500970 480 502250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 500970 709904 502250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 508970 480 510250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 508970 709904 510250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 516970 480 518250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 516970 709904 518250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 524970 480 526250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 524970 709904 526250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 532970 480 534250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 532970 709904 534250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 540970 480 542250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 540970 709904 542250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 548970 480 550250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 548970 709904 550250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 556970 480 558250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 556970 709904 558250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 564970 480 566250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 564970 709904 566250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 572970 480 574250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 572970 709904 574250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 580970 480 582250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 580970 709904 582250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 588970 480 590250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 588970 709904 590250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 596970 480 598250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 596970 709904 598250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 604970 480 606250 389968 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 604970 709904 606250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 612970 480 614250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 620970 480 622250 952608 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 14006 633004 15286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 22006 633004 23286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 30006 633004 31286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 38006 633004 39286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 46006 633004 47286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 54006 633004 55286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 62006 633004 63286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 70006 633004 71286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 78006 633004 79286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 86006 633004 87286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 94006 633004 95286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 102006 633004 103286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 110006 633004 111286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 118006 633004 119286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 126006 633004 127286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 134006 633004 135286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 142006 633004 143286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 150006 633004 151286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 158006 633004 159286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 166006 633004 167286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 174006 633004 175286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 182006 633004 183286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 190006 633004 191286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 198006 633004 199286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 206006 633004 207286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 214006 633004 215286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 222006 633004 223286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 230006 633004 231286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 238006 633004 239286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 246006 633004 247286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 254006 633004 255286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 262006 633004 263286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 270006 633004 271286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 278006 633004 279286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 286006 633004 287286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 294006 633004 295286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 302006 633004 303286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 310006 633004 311286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 318006 633004 319286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 326006 633004 327286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 334006 633004 335286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 342006 633004 343286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 350006 633004 351286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 358006 633004 359286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 366006 633004 367286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 374006 633004 375286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 382006 633004 383286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 390006 633004 391286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 398006 633004 399286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 406006 633004 407286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 414006 633004 415286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 422006 633004 423286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 430006 633004 431286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 438006 633004 439286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 446006 633004 447286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 454006 139548 455286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 462006 139548 463286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 470006 139548 471286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 478006 139548 479286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 486006 139548 487286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 494006 139548 495286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 502006 139548 503286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 510006 139548 511286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 518006 139548 519286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 526006 139548 527286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 534006 139548 535286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 542006 139548 543286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 550006 633004 551286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 558006 633004 559286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 566006 633004 567286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 574006 633004 575286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 582006 633004 583286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 590006 633004 591286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 598006 633004 599286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 606006 633004 607286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 614006 633004 615286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 622006 633004 623286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 630006 633004 631286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 638006 633004 639286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 646006 633004 647286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 654006 633004 655286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 662006 633004 663286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 670006 633004 671286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 678006 633004 679286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 686006 633004 687286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 694006 633004 695286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 702006 633004 703286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 710006 633004 711286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 718006 633004 719286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 726006 633004 727286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 734006 633004 735286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 742006 633004 743286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 750006 633004 751286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 758006 633004 759286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 766006 633004 767286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 774006 633004 775286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 782006 633004 783286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 790006 633004 791286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 798006 633004 799286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 806006 633004 807286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 814006 633004 815286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 822006 633004 823286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 830006 633004 831286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 838006 633004 839286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 846006 633004 847286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 854006 633004 855286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 862006 633004 863286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 870006 633004 871286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 878006 633004 879286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 886006 633004 887286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 894006 633004 895286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 902006 633004 903286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 910006 633004 911286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 918006 633004 919286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 926006 633004 927286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 934006 633004 935286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 324 942006 633004 943286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 454006 633004 455286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 462006 633004 463286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 470006 633004 471286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 478006 633004 479286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 486006 633004 487286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 494006 633004 495286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 502006 633004 503286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 510006 633004 511286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 518006 633004 519286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 526006 633004 527286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 534006 633004 535286 6 vssd1
port 875 nsew ground bidirectional
rlabel metal5 s 433660 542006 633004 543286 6 vssd1
port 875 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 633326 953326
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 666563062
string GDS_FILE /home/hosni/caravel_openframe_project/openlane/openframe_project_wrapper/runs/23_09_17_16_29/results/signoff/openframe_project_wrapper.magic.gds
string GDS_START 220471022
<< end >>

