VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO picosoc
  CLASS BLOCK ;
  FOREIGN picosoc ;
  ORIGIN 0.000 0.000 ;
  SIZE 2600.000 BY 1600.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.070 10.640 17.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 10.640 57.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.070 10.640 97.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.070 1046.620 97.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.070 10.640 137.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.070 1046.620 137.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.070 10.640 177.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.070 1046.620 177.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.070 10.640 217.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.070 1046.620 217.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.070 10.640 257.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.070 1047.240 257.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.070 10.640 297.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.070 1046.620 297.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.070 10.640 337.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.070 1046.620 337.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.070 10.640 377.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.070 1046.620 377.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.070 10.640 417.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.070 1046.620 417.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.070 10.640 457.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.070 1047.240 457.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.070 10.640 497.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.070 1046.620 497.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.070 10.640 537.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.070 1046.620 537.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.070 10.640 577.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.070 1046.620 577.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.070 10.640 617.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 614.070 1047.240 617.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.070 10.640 657.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.070 1046.620 657.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.070 10.640 697.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.070 1046.620 697.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 734.070 10.640 737.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 734.070 1046.620 737.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.070 10.640 777.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.070 1046.620 777.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.070 10.640 817.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.070 10.640 857.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.070 10.640 897.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 934.070 10.640 937.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.070 10.640 977.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1014.070 10.640 1017.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.070 10.640 1057.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1094.070 10.640 1097.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1134.070 10.640 1137.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1174.070 10.640 1177.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.070 10.640 1217.170 741.155 ;
    END
    PORT
      LAYER met4 ;
        RECT 1214.070 770.365 1217.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.070 10.640 1257.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1294.070 10.640 1297.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1334.070 10.640 1337.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.070 10.640 1377.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.070 10.640 1417.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.070 1046.620 1417.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.070 10.640 1457.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.070 1046.620 1457.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1494.070 10.640 1497.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1494.070 1046.620 1497.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.070 10.640 1537.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1534.070 1046.620 1537.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1574.070 10.640 1577.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1574.070 1046.620 1577.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.070 10.640 1617.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1614.070 1047.240 1617.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.070 10.640 1657.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.070 1047.240 1657.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1694.070 10.640 1697.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1694.070 1046.620 1697.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1734.070 10.640 1737.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1734.070 1046.620 1737.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.070 10.640 1777.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.070 1046.620 1777.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.070 10.640 1817.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1814.070 1047.240 1817.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.070 10.640 1857.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.070 1047.240 1857.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.070 10.640 1897.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.070 1046.620 1897.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.070 10.640 1937.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1934.070 1046.620 1937.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1974.070 10.640 1977.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1974.070 1046.620 1977.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2014.070 10.640 2017.170 609.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2014.070 1046.620 2017.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.070 10.640 2057.170 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.070 1047.240 2057.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.070 10.640 2097.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.070 10.640 2137.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.070 10.640 2177.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2214.070 10.640 2217.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.070 10.640 2257.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2294.070 10.640 2297.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2334.070 10.640 2337.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.070 10.640 2377.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2414.070 10.640 2417.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.070 10.640 2457.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.070 10.640 2497.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2534.070 10.640 2537.170 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2574.070 10.640 2577.170 1588.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.430 2594.640 22.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 59.430 2594.640 62.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 99.430 2594.640 102.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 139.430 2594.640 142.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.430 2594.640 182.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 219.430 2594.640 222.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 259.430 2594.640 262.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 299.430 2594.640 302.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 339.430 2594.640 342.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 379.430 2594.640 382.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 419.430 2594.640 422.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 459.430 2594.640 462.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 499.430 2594.640 502.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 539.430 2594.640 542.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 579.430 2594.640 582.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 619.430 2594.640 622.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 659.430 2594.640 662.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 699.430 2594.640 702.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 739.430 2594.640 742.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 779.430 2594.640 782.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 819.430 2594.640 822.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 859.430 2594.640 862.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 899.430 2594.640 902.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 939.430 2594.640 942.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 979.430 2594.640 982.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1019.430 2594.640 1022.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1059.430 2594.640 1062.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1099.430 2594.640 1102.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1139.430 2594.640 1142.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1179.430 2594.640 1182.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1219.430 2594.640 1222.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1259.430 2594.640 1262.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1299.430 2594.640 1302.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1339.430 2594.640 1342.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1379.430 2594.640 1382.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1419.430 2594.640 1422.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1459.430 2594.640 1462.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1499.430 2594.640 1502.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1539.430 2594.640 1542.530 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1579.430 2594.640 1582.530 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.970 10.640 52.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.970 10.640 92.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.970 1046.620 92.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.970 10.640 132.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 128.970 1046.620 132.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.970 10.640 172.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.970 1046.620 172.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 10.640 212.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.970 1046.620 212.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.970 10.640 252.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.970 1046.620 252.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 10.640 292.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.970 1046.960 292.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.970 10.640 332.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.970 1046.960 332.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1046.620 372.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 10.640 412.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.970 1046.620 412.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.970 10.640 452.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.970 1046.620 452.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.970 10.640 492.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 488.970 1046.620 492.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 528.970 10.640 532.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 528.970 1046.960 532.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 10.640 572.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.970 1046.620 572.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 10.640 612.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.970 1046.620 612.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.970 10.640 652.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 648.970 1046.620 652.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 688.970 10.640 692.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 688.970 1046.960 692.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1046.620 732.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 768.970 10.640 772.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 768.970 1046.620 772.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.970 10.640 812.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 848.970 10.640 852.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 888.970 10.640 892.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 928.970 10.640 932.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 968.970 10.640 972.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.970 10.640 1012.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1048.970 10.640 1052.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1128.970 10.640 1132.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1168.970 10.640 1172.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 10.640 1212.070 694.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.970 778.940 1212.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1248.970 10.640 1252.070 694.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1248.970 778.940 1252.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1288.970 10.640 1292.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1328.970 10.640 1332.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1368.970 10.640 1372.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 10.640 1412.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.970 1046.620 1412.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 10.640 1452.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 1046.620 1452.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1488.970 10.640 1492.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1488.970 1046.620 1492.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1528.970 10.640 1532.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1528.970 1046.620 1532.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1568.970 10.640 1572.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1568.970 1046.620 1572.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 10.640 1612.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.970 1046.620 1612.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1648.970 10.640 1652.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1648.970 1046.620 1652.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 10.640 1692.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1688.970 1046.960 1692.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.970 10.640 1732.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1728.970 1046.960 1732.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.970 10.640 1772.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1768.970 1046.620 1772.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 10.640 1812.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1046.620 1812.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.970 10.640 1852.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1848.970 1046.620 1852.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1888.970 10.640 1892.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1888.970 1046.960 1892.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1928.970 10.640 1932.070 609.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1928.970 1046.960 1932.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 10.640 1972.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1968.970 1046.620 1972.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 10.640 2012.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 1046.620 2012.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.970 10.640 2052.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2048.970 1046.620 2052.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2088.970 10.640 2092.070 609.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2088.970 1046.620 2092.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2128.970 10.640 2132.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 10.640 2172.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.970 10.640 2212.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.970 10.640 2252.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2288.970 10.640 2292.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2328.970 10.640 2332.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2368.970 10.640 2372.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.970 10.640 2412.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2448.970 10.640 2452.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2488.970 10.640 2492.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 10.640 2532.070 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2568.970 10.640 2572.070 1588.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.330 2594.640 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 54.330 2594.640 57.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 94.330 2594.640 97.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 134.330 2594.640 137.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 174.330 2594.640 177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 214.330 2594.640 217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 254.330 2594.640 257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 294.330 2594.640 297.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 334.330 2594.640 337.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 374.330 2594.640 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 414.330 2594.640 417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 454.330 2594.640 457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 494.330 2594.640 497.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 534.330 2594.640 537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 574.330 2594.640 577.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 614.330 2594.640 617.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 654.330 2594.640 657.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 694.330 2594.640 697.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 734.330 2594.640 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 774.330 2594.640 777.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 814.330 2594.640 817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 854.330 2594.640 857.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 894.330 2594.640 897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 934.330 2594.640 937.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 974.330 2594.640 977.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1014.330 2594.640 1017.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1054.330 2594.640 1057.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1094.330 2594.640 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1134.330 2594.640 1137.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1174.330 2594.640 1177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1214.330 2594.640 1217.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1254.330 2594.640 1257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1294.330 2594.640 1297.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1334.330 2594.640 1337.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1374.330 2594.640 1377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1414.330 2594.640 1417.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1454.330 2594.640 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1494.330 2594.640 1497.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1534.330 2594.640 1537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1574.330 2594.640 1577.430 ;
    END
  END VPWR
  PIN gpio_dm0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 93.880 2600.000 94.480 ;
    END
  END gpio_dm0[0]
  PIN gpio_dm0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1073.080 2600.000 1073.680 ;
    END
  END gpio_dm0[10]
  PIN gpio_dm0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1171.000 2600.000 1171.600 ;
    END
  END gpio_dm0[11]
  PIN gpio_dm0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1268.920 2600.000 1269.520 ;
    END
  END gpio_dm0[12]
  PIN gpio_dm0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1366.840 2600.000 1367.440 ;
    END
  END gpio_dm0[13]
  PIN gpio_dm0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1464.760 2600.000 1465.360 ;
    END
  END gpio_dm0[14]
  PIN gpio_dm0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2507.550 1597.600 2507.830 1600.000 ;
    END
  END gpio_dm0[15]
  PIN gpio_dm0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2220.510 1597.600 2220.790 1600.000 ;
    END
  END gpio_dm0[16]
  PIN gpio_dm0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1933.470 1597.600 1933.750 1600.000 ;
    END
  END gpio_dm0[17]
  PIN gpio_dm0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1646.430 1597.600 1646.710 1600.000 ;
    END
  END gpio_dm0[18]
  PIN gpio_dm0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1359.390 1597.600 1359.670 1600.000 ;
    END
  END gpio_dm0[19]
  PIN gpio_dm0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 191.800 2600.000 192.400 ;
    END
  END gpio_dm0[1]
  PIN gpio_dm0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1597.600 1072.630 1600.000 ;
    END
  END gpio_dm0[20]
  PIN gpio_dm0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 785.310 1597.600 785.590 1600.000 ;
    END
  END gpio_dm0[21]
  PIN gpio_dm0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 498.270 1597.600 498.550 1600.000 ;
    END
  END gpio_dm0[22]
  PIN gpio_dm0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 211.230 1597.600 211.510 1600.000 ;
    END
  END gpio_dm0[23]
  PIN gpio_dm0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1464.760 2.400 1465.360 ;
    END
  END gpio_dm0[24]
  PIN gpio_dm0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 2.400 1367.440 ;
    END
  END gpio_dm0[25]
  PIN gpio_dm0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.920 2.400 1269.520 ;
    END
  END gpio_dm0[26]
  PIN gpio_dm0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1171.000 2.400 1171.600 ;
    END
  END gpio_dm0[27]
  PIN gpio_dm0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.080 2.400 1073.680 ;
    END
  END gpio_dm0[28]
  PIN gpio_dm0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 2.400 975.760 ;
    END
  END gpio_dm0[29]
  PIN gpio_dm0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 289.720 2600.000 290.320 ;
    END
  END gpio_dm0[2]
  PIN gpio_dm0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 2.400 877.840 ;
    END
  END gpio_dm0[30]
  PIN gpio_dm0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 2.400 779.920 ;
    END
  END gpio_dm0[31]
  PIN gpio_dm0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 2.400 682.000 ;
    END
  END gpio_dm0[32]
  PIN gpio_dm0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 2.400 584.080 ;
    END
  END gpio_dm0[33]
  PIN gpio_dm0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 2.400 486.160 ;
    END
  END gpio_dm0[34]
  PIN gpio_dm0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 2.400 388.240 ;
    END
  END gpio_dm0[35]
  PIN gpio_dm0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 2.400 290.320 ;
    END
  END gpio_dm0[36]
  PIN gpio_dm0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 2.400 192.400 ;
    END
  END gpio_dm0[37]
  PIN gpio_dm0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 2.400 ;
    END
  END gpio_dm0[38]
  PIN gpio_dm0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 2.400 ;
    END
  END gpio_dm0[39]
  PIN gpio_dm0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 387.640 2600.000 388.240 ;
    END
  END gpio_dm0[3]
  PIN gpio_dm0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 2.400 ;
    END
  END gpio_dm0[40]
  PIN gpio_dm0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1007.030 0.000 1007.310 2.400 ;
    END
  END gpio_dm0[41]
  PIN gpio_dm0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 2.400 ;
    END
  END gpio_dm0[42]
  PIN gpio_dm0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1592.150 0.000 1592.430 2.400 ;
    END
  END gpio_dm0[43]
  PIN gpio_dm0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 485.560 2600.000 486.160 ;
    END
  END gpio_dm0[4]
  PIN gpio_dm0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 583.480 2600.000 584.080 ;
    END
  END gpio_dm0[5]
  PIN gpio_dm0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 681.400 2600.000 682.000 ;
    END
  END gpio_dm0[6]
  PIN gpio_dm0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 779.320 2600.000 779.920 ;
    END
  END gpio_dm0[7]
  PIN gpio_dm0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 877.240 2600.000 877.840 ;
    END
  END gpio_dm0[8]
  PIN gpio_dm0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 975.160 2600.000 975.760 ;
    END
  END gpio_dm0[9]
  PIN gpio_dm1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 85.720 2600.000 86.320 ;
    END
  END gpio_dm1[0]
  PIN gpio_dm1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1064.920 2600.000 1065.520 ;
    END
  END gpio_dm1[10]
  PIN gpio_dm1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1162.840 2600.000 1163.440 ;
    END
  END gpio_dm1[11]
  PIN gpio_dm1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1260.760 2600.000 1261.360 ;
    END
  END gpio_dm1[12]
  PIN gpio_dm1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1358.680 2600.000 1359.280 ;
    END
  END gpio_dm1[13]
  PIN gpio_dm1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1456.600 2600.000 1457.200 ;
    END
  END gpio_dm1[14]
  PIN gpio_dm1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2531.470 1597.600 2531.750 1600.000 ;
    END
  END gpio_dm1[15]
  PIN gpio_dm1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2244.430 1597.600 2244.710 1600.000 ;
    END
  END gpio_dm1[16]
  PIN gpio_dm1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1957.390 1597.600 1957.670 1600.000 ;
    END
  END gpio_dm1[17]
  PIN gpio_dm1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1670.350 1597.600 1670.630 1600.000 ;
    END
  END gpio_dm1[18]
  PIN gpio_dm1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1383.310 1597.600 1383.590 1600.000 ;
    END
  END gpio_dm1[19]
  PIN gpio_dm1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 183.640 2600.000 184.240 ;
    END
  END gpio_dm1[1]
  PIN gpio_dm1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1096.270 1597.600 1096.550 1600.000 ;
    END
  END gpio_dm1[20]
  PIN gpio_dm1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 809.230 1597.600 809.510 1600.000 ;
    END
  END gpio_dm1[21]
  PIN gpio_dm1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 522.190 1597.600 522.470 1600.000 ;
    END
  END gpio_dm1[22]
  PIN gpio_dm1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 235.150 1597.600 235.430 1600.000 ;
    END
  END gpio_dm1[23]
  PIN gpio_dm1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 2.400 1473.520 ;
    END
  END gpio_dm1[24]
  PIN gpio_dm1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.000 2.400 1375.600 ;
    END
  END gpio_dm1[25]
  PIN gpio_dm1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.080 2.400 1277.680 ;
    END
  END gpio_dm1[26]
  PIN gpio_dm1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.160 2.400 1179.760 ;
    END
  END gpio_dm1[27]
  PIN gpio_dm1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 2.400 1081.840 ;
    END
  END gpio_dm1[28]
  PIN gpio_dm1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 2.400 983.920 ;
    END
  END gpio_dm1[29]
  PIN gpio_dm1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 281.560 2600.000 282.160 ;
    END
  END gpio_dm1[2]
  PIN gpio_dm1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.400 2.400 886.000 ;
    END
  END gpio_dm1[30]
  PIN gpio_dm1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 2.400 788.080 ;
    END
  END gpio_dm1[31]
  PIN gpio_dm1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 2.400 690.160 ;
    END
  END gpio_dm1[32]
  PIN gpio_dm1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 2.400 592.240 ;
    END
  END gpio_dm1[33]
  PIN gpio_dm1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 2.400 494.320 ;
    END
  END gpio_dm1[34]
  PIN gpio_dm1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 2.400 396.400 ;
    END
  END gpio_dm1[35]
  PIN gpio_dm1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 2.400 298.480 ;
    END
  END gpio_dm1[36]
  PIN gpio_dm1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 2.400 200.560 ;
    END
  END gpio_dm1[37]
  PIN gpio_dm1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END gpio_dm1[38]
  PIN gpio_dm1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 2.400 ;
    END
  END gpio_dm1[39]
  PIN gpio_dm1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 379.480 2600.000 380.080 ;
    END
  END gpio_dm1[3]
  PIN gpio_dm1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 2.400 ;
    END
  END gpio_dm1[40]
  PIN gpio_dm1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 982.650 0.000 982.930 2.400 ;
    END
  END gpio_dm1[41]
  PIN gpio_dm1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1275.210 0.000 1275.490 2.400 ;
    END
  END gpio_dm1[42]
  PIN gpio_dm1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1567.770 0.000 1568.050 2.400 ;
    END
  END gpio_dm1[43]
  PIN gpio_dm1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 477.400 2600.000 478.000 ;
    END
  END gpio_dm1[4]
  PIN gpio_dm1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 575.320 2600.000 575.920 ;
    END
  END gpio_dm1[5]
  PIN gpio_dm1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 673.240 2600.000 673.840 ;
    END
  END gpio_dm1[6]
  PIN gpio_dm1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 771.160 2600.000 771.760 ;
    END
  END gpio_dm1[7]
  PIN gpio_dm1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 869.080 2600.000 869.680 ;
    END
  END gpio_dm1[8]
  PIN gpio_dm1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 967.000 2600.000 967.600 ;
    END
  END gpio_dm1[9]
  PIN gpio_dm2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 110.200 2600.000 110.800 ;
    END
  END gpio_dm2[0]
  PIN gpio_dm2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1089.400 2600.000 1090.000 ;
    END
  END gpio_dm2[10]
  PIN gpio_dm2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1187.320 2600.000 1187.920 ;
    END
  END gpio_dm2[11]
  PIN gpio_dm2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1285.240 2600.000 1285.840 ;
    END
  END gpio_dm2[12]
  PIN gpio_dm2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1383.160 2600.000 1383.760 ;
    END
  END gpio_dm2[13]
  PIN gpio_dm2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1481.080 2600.000 1481.680 ;
    END
  END gpio_dm2[14]
  PIN gpio_dm2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2459.710 1597.600 2459.990 1600.000 ;
    END
  END gpio_dm2[15]
  PIN gpio_dm2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2172.670 1597.600 2172.950 1600.000 ;
    END
  END gpio_dm2[16]
  PIN gpio_dm2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1885.630 1597.600 1885.910 1600.000 ;
    END
  END gpio_dm2[17]
  PIN gpio_dm2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1598.590 1597.600 1598.870 1600.000 ;
    END
  END gpio_dm2[18]
  PIN gpio_dm2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1311.550 1597.600 1311.830 1600.000 ;
    END
  END gpio_dm2[19]
  PIN gpio_dm2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 208.120 2600.000 208.720 ;
    END
  END gpio_dm2[1]
  PIN gpio_dm2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1024.510 1597.600 1024.790 1600.000 ;
    END
  END gpio_dm2[20]
  PIN gpio_dm2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 737.470 1597.600 737.750 1600.000 ;
    END
  END gpio_dm2[21]
  PIN gpio_dm2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 450.430 1597.600 450.710 1600.000 ;
    END
  END gpio_dm2[22]
  PIN gpio_dm2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 163.390 1597.600 163.670 1600.000 ;
    END
  END gpio_dm2[23]
  PIN gpio_dm2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 2.400 1449.040 ;
    END
  END gpio_dm2[24]
  PIN gpio_dm2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1350.520 2.400 1351.120 ;
    END
  END gpio_dm2[25]
  PIN gpio_dm2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1252.600 2.400 1253.200 ;
    END
  END gpio_dm2[26]
  PIN gpio_dm2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.680 2.400 1155.280 ;
    END
  END gpio_dm2[27]
  PIN gpio_dm2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.760 2.400 1057.360 ;
    END
  END gpio_dm2[28]
  PIN gpio_dm2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 2.400 959.440 ;
    END
  END gpio_dm2[29]
  PIN gpio_dm2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 306.040 2600.000 306.640 ;
    END
  END gpio_dm2[2]
  PIN gpio_dm2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 2.400 861.520 ;
    END
  END gpio_dm2[30]
  PIN gpio_dm2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 2.400 763.600 ;
    END
  END gpio_dm2[31]
  PIN gpio_dm2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 2.400 665.680 ;
    END
  END gpio_dm2[32]
  PIN gpio_dm2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 2.400 567.760 ;
    END
  END gpio_dm2[33]
  PIN gpio_dm2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 2.400 469.840 ;
    END
  END gpio_dm2[34]
  PIN gpio_dm2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 2.400 371.920 ;
    END
  END gpio_dm2[35]
  PIN gpio_dm2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 2.400 274.000 ;
    END
  END gpio_dm2[36]
  PIN gpio_dm2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 2.400 176.080 ;
    END
  END gpio_dm2[37]
  PIN gpio_dm2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 2.400 ;
    END
  END gpio_dm2[38]
  PIN gpio_dm2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 2.400 ;
    END
  END gpio_dm2[39]
  PIN gpio_dm2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 403.960 2600.000 404.560 ;
    END
  END gpio_dm2[3]
  PIN gpio_dm2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 2.400 ;
    END
  END gpio_dm2[40]
  PIN gpio_dm2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 2.400 ;
    END
  END gpio_dm2[41]
  PIN gpio_dm2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 2.400 ;
    END
  END gpio_dm2[42]
  PIN gpio_dm2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1640.910 0.000 1641.190 2.400 ;
    END
  END gpio_dm2[43]
  PIN gpio_dm2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 501.880 2600.000 502.480 ;
    END
  END gpio_dm2[4]
  PIN gpio_dm2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 599.800 2600.000 600.400 ;
    END
  END gpio_dm2[5]
  PIN gpio_dm2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 697.720 2600.000 698.320 ;
    END
  END gpio_dm2[6]
  PIN gpio_dm2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 795.640 2600.000 796.240 ;
    END
  END gpio_dm2[7]
  PIN gpio_dm2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 893.560 2600.000 894.160 ;
    END
  END gpio_dm2[8]
  PIN gpio_dm2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 991.480 2600.000 992.080 ;
    END
  END gpio_dm2[9]
  PIN gpio_ib_mode_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 134.680 2600.000 135.280 ;
    END
  END gpio_ib_mode_sel[0]
  PIN gpio_ib_mode_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1113.880 2600.000 1114.480 ;
    END
  END gpio_ib_mode_sel[10]
  PIN gpio_ib_mode_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1211.800 2600.000 1212.400 ;
    END
  END gpio_ib_mode_sel[11]
  PIN gpio_ib_mode_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1309.720 2600.000 1310.320 ;
    END
  END gpio_ib_mode_sel[12]
  PIN gpio_ib_mode_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1407.640 2600.000 1408.240 ;
    END
  END gpio_ib_mode_sel[13]
  PIN gpio_ib_mode_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1505.560 2600.000 1506.160 ;
    END
  END gpio_ib_mode_sel[14]
  PIN gpio_ib_mode_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2387.950 1597.600 2388.230 1600.000 ;
    END
  END gpio_ib_mode_sel[15]
  PIN gpio_ib_mode_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2100.910 1597.600 2101.190 1600.000 ;
    END
  END gpio_ib_mode_sel[16]
  PIN gpio_ib_mode_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1813.870 1597.600 1814.150 1600.000 ;
    END
  END gpio_ib_mode_sel[17]
  PIN gpio_ib_mode_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1526.830 1597.600 1527.110 1600.000 ;
    END
  END gpio_ib_mode_sel[18]
  PIN gpio_ib_mode_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1239.790 1597.600 1240.070 1600.000 ;
    END
  END gpio_ib_mode_sel[19]
  PIN gpio_ib_mode_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 232.600 2600.000 233.200 ;
    END
  END gpio_ib_mode_sel[1]
  PIN gpio_ib_mode_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 952.750 1597.600 953.030 1600.000 ;
    END
  END gpio_ib_mode_sel[20]
  PIN gpio_ib_mode_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 665.710 1597.600 665.990 1600.000 ;
    END
  END gpio_ib_mode_sel[21]
  PIN gpio_ib_mode_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 378.670 1597.600 378.950 1600.000 ;
    END
  END gpio_ib_mode_sel[22]
  PIN gpio_ib_mode_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 91.630 1597.600 91.910 1600.000 ;
    END
  END gpio_ib_mode_sel[23]
  PIN gpio_ib_mode_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.960 2.400 1424.560 ;
    END
  END gpio_ib_mode_sel[24]
  PIN gpio_ib_mode_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 2.400 1326.640 ;
    END
  END gpio_ib_mode_sel[25]
  PIN gpio_ib_mode_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1228.120 2.400 1228.720 ;
    END
  END gpio_ib_mode_sel[26]
  PIN gpio_ib_mode_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.200 2.400 1130.800 ;
    END
  END gpio_ib_mode_sel[27]
  PIN gpio_ib_mode_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 2.400 1032.880 ;
    END
  END gpio_ib_mode_sel[28]
  PIN gpio_ib_mode_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 2.400 934.960 ;
    END
  END gpio_ib_mode_sel[29]
  PIN gpio_ib_mode_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 330.520 2600.000 331.120 ;
    END
  END gpio_ib_mode_sel[2]
  PIN gpio_ib_mode_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 2.400 837.040 ;
    END
  END gpio_ib_mode_sel[30]
  PIN gpio_ib_mode_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 2.400 739.120 ;
    END
  END gpio_ib_mode_sel[31]
  PIN gpio_ib_mode_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 2.400 641.200 ;
    END
  END gpio_ib_mode_sel[32]
  PIN gpio_ib_mode_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 2.400 543.280 ;
    END
  END gpio_ib_mode_sel[33]
  PIN gpio_ib_mode_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 2.400 445.360 ;
    END
  END gpio_ib_mode_sel[34]
  PIN gpio_ib_mode_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 2.400 347.440 ;
    END
  END gpio_ib_mode_sel[35]
  PIN gpio_ib_mode_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 2.400 249.520 ;
    END
  END gpio_ib_mode_sel[36]
  PIN gpio_ib_mode_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 2.400 151.600 ;
    END
  END gpio_ib_mode_sel[37]
  PIN gpio_ib_mode_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 2.400 ;
    END
  END gpio_ib_mode_sel[38]
  PIN gpio_ib_mode_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 2.400 ;
    END
  END gpio_ib_mode_sel[39]
  PIN gpio_ib_mode_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 428.440 2600.000 429.040 ;
    END
  END gpio_ib_mode_sel[3]
  PIN gpio_ib_mode_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 2.400 ;
    END
  END gpio_ib_mode_sel[40]
  PIN gpio_ib_mode_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 2.400 ;
    END
  END gpio_ib_mode_sel[41]
  PIN gpio_ib_mode_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1421.490 0.000 1421.770 2.400 ;
    END
  END gpio_ib_mode_sel[42]
  PIN gpio_ib_mode_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1714.050 0.000 1714.330 2.400 ;
    END
  END gpio_ib_mode_sel[43]
  PIN gpio_ib_mode_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 526.360 2600.000 526.960 ;
    END
  END gpio_ib_mode_sel[4]
  PIN gpio_ib_mode_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 624.280 2600.000 624.880 ;
    END
  END gpio_ib_mode_sel[5]
  PIN gpio_ib_mode_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 722.200 2600.000 722.800 ;
    END
  END gpio_ib_mode_sel[6]
  PIN gpio_ib_mode_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 820.120 2600.000 820.720 ;
    END
  END gpio_ib_mode_sel[7]
  PIN gpio_ib_mode_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 918.040 2600.000 918.640 ;
    END
  END gpio_ib_mode_sel[8]
  PIN gpio_ib_mode_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1015.960 2600.000 1016.560 ;
    END
  END gpio_ib_mode_sel[9]
  PIN gpio_ieb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 102.040 2600.000 102.640 ;
    END
  END gpio_ieb[0]
  PIN gpio_ieb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1081.240 2600.000 1081.840 ;
    END
  END gpio_ieb[10]
  PIN gpio_ieb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1179.160 2600.000 1179.760 ;
    END
  END gpio_ieb[11]
  PIN gpio_ieb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1277.080 2600.000 1277.680 ;
    END
  END gpio_ieb[12]
  PIN gpio_ieb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1375.000 2600.000 1375.600 ;
    END
  END gpio_ieb[13]
  PIN gpio_ieb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1472.920 2600.000 1473.520 ;
    END
  END gpio_ieb[14]
  PIN gpio_ieb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2483.630 1597.600 2483.910 1600.000 ;
    END
  END gpio_ieb[15]
  PIN gpio_ieb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2196.590 1597.600 2196.870 1600.000 ;
    END
  END gpio_ieb[16]
  PIN gpio_ieb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1909.550 1597.600 1909.830 1600.000 ;
    END
  END gpio_ieb[17]
  PIN gpio_ieb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1622.510 1597.600 1622.790 1600.000 ;
    END
  END gpio_ieb[18]
  PIN gpio_ieb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1335.470 1597.600 1335.750 1600.000 ;
    END
  END gpio_ieb[19]
  PIN gpio_ieb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 199.960 2600.000 200.560 ;
    END
  END gpio_ieb[1]
  PIN gpio_ieb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1048.430 1597.600 1048.710 1600.000 ;
    END
  END gpio_ieb[20]
  PIN gpio_ieb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 761.390 1597.600 761.670 1600.000 ;
    END
  END gpio_ieb[21]
  PIN gpio_ieb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 474.350 1597.600 474.630 1600.000 ;
    END
  END gpio_ieb[22]
  PIN gpio_ieb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 187.310 1597.600 187.590 1600.000 ;
    END
  END gpio_ieb[23]
  PIN gpio_ieb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1456.600 2.400 1457.200 ;
    END
  END gpio_ieb[24]
  PIN gpio_ieb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1358.680 2.400 1359.280 ;
    END
  END gpio_ieb[25]
  PIN gpio_ieb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 2.400 1261.360 ;
    END
  END gpio_ieb[26]
  PIN gpio_ieb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 2.400 1163.440 ;
    END
  END gpio_ieb[27]
  PIN gpio_ieb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 2.400 1065.520 ;
    END
  END gpio_ieb[28]
  PIN gpio_ieb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.000 2.400 967.600 ;
    END
  END gpio_ieb[29]
  PIN gpio_ieb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 297.880 2600.000 298.480 ;
    END
  END gpio_ieb[2]
  PIN gpio_ieb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.080 2.400 869.680 ;
    END
  END gpio_ieb[30]
  PIN gpio_ieb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 2.400 771.760 ;
    END
  END gpio_ieb[31]
  PIN gpio_ieb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 2.400 673.840 ;
    END
  END gpio_ieb[32]
  PIN gpio_ieb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 2.400 575.920 ;
    END
  END gpio_ieb[33]
  PIN gpio_ieb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 2.400 478.000 ;
    END
  END gpio_ieb[34]
  PIN gpio_ieb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 2.400 380.080 ;
    END
  END gpio_ieb[35]
  PIN gpio_ieb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 2.400 282.160 ;
    END
  END gpio_ieb[36]
  PIN gpio_ieb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 2.400 184.240 ;
    END
  END gpio_ieb[37]
  PIN gpio_ieb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 2.400 ;
    END
  END gpio_ieb[38]
  PIN gpio_ieb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 2.400 ;
    END
  END gpio_ieb[39]
  PIN gpio_ieb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 395.800 2600.000 396.400 ;
    END
  END gpio_ieb[3]
  PIN gpio_ieb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 2.400 ;
    END
  END gpio_ieb[40]
  PIN gpio_ieb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1031.410 0.000 1031.690 2.400 ;
    END
  END gpio_ieb[41]
  PIN gpio_ieb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 2.400 ;
    END
  END gpio_ieb[42]
  PIN gpio_ieb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1616.530 0.000 1616.810 2.400 ;
    END
  END gpio_ieb[43]
  PIN gpio_ieb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 493.720 2600.000 494.320 ;
    END
  END gpio_ieb[4]
  PIN gpio_ieb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 591.640 2600.000 592.240 ;
    END
  END gpio_ieb[5]
  PIN gpio_ieb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 689.560 2600.000 690.160 ;
    END
  END gpio_ieb[6]
  PIN gpio_ieb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 787.480 2600.000 788.080 ;
    END
  END gpio_ieb[7]
  PIN gpio_ieb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 885.400 2600.000 886.000 ;
    END
  END gpio_ieb[8]
  PIN gpio_ieb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 983.320 2600.000 983.920 ;
    END
  END gpio_ieb[9]
  PIN gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 69.400 2600.000 70.000 ;
    END
  END gpio_in[0]
  PIN gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1048.600 2600.000 1049.200 ;
    END
  END gpio_in[10]
  PIN gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1146.520 2600.000 1147.120 ;
    END
  END gpio_in[11]
  PIN gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1244.440 2600.000 1245.040 ;
    END
  END gpio_in[12]
  PIN gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1342.360 2600.000 1342.960 ;
    END
  END gpio_in[13]
  PIN gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1440.280 2600.000 1440.880 ;
    END
  END gpio_in[14]
  PIN gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2579.310 1597.600 2579.590 1600.000 ;
    END
  END gpio_in[15]
  PIN gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2292.270 1597.600 2292.550 1600.000 ;
    END
  END gpio_in[16]
  PIN gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2005.230 1597.600 2005.510 1600.000 ;
    END
  END gpio_in[17]
  PIN gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1718.190 1597.600 1718.470 1600.000 ;
    END
  END gpio_in[18]
  PIN gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1431.150 1597.600 1431.430 1600.000 ;
    END
  END gpio_in[19]
  PIN gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 167.320 2600.000 167.920 ;
    END
  END gpio_in[1]
  PIN gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1144.110 1597.600 1144.390 1600.000 ;
    END
  END gpio_in[20]
  PIN gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 857.070 1597.600 857.350 1600.000 ;
    END
  END gpio_in[21]
  PIN gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 570.030 1597.600 570.310 1600.000 ;
    END
  END gpio_in[22]
  PIN gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 282.990 1597.600 283.270 1600.000 ;
    END
  END gpio_in[23]
  PIN gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 2.400 1489.840 ;
    END
  END gpio_in[24]
  PIN gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1391.320 2.400 1391.920 ;
    END
  END gpio_in[25]
  PIN gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 2.400 1294.000 ;
    END
  END gpio_in[26]
  PIN gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1195.480 2.400 1196.080 ;
    END
  END gpio_in[27]
  PIN gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1097.560 2.400 1098.160 ;
    END
  END gpio_in[28]
  PIN gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 2.400 1000.240 ;
    END
  END gpio_in[29]
  PIN gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 265.240 2600.000 265.840 ;
    END
  END gpio_in[2]
  PIN gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 2.400 902.320 ;
    END
  END gpio_in[30]
  PIN gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 2.400 804.400 ;
    END
  END gpio_in[31]
  PIN gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 2.400 706.480 ;
    END
  END gpio_in[32]
  PIN gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 2.400 608.560 ;
    END
  END gpio_in[33]
  PIN gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 2.400 510.640 ;
    END
  END gpio_in[34]
  PIN gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 2.400 412.720 ;
    END
  END gpio_in[35]
  PIN gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 2.400 314.800 ;
    END
  END gpio_in[36]
  PIN gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 2.400 216.880 ;
    END
  END gpio_in[37]
  PIN gpio_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END gpio_in[38]
  PIN gpio_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 2.400 ;
    END
  END gpio_in[39]
  PIN gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 363.160 2600.000 363.760 ;
    END
  END gpio_in[3]
  PIN gpio_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 2.400 ;
    END
  END gpio_in[40]
  PIN gpio_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 2.400 ;
    END
  END gpio_in[41]
  PIN gpio_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 2.400 ;
    END
  END gpio_in[42]
  PIN gpio_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1519.010 0.000 1519.290 2.400 ;
    END
  END gpio_in[43]
  PIN gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 461.080 2600.000 461.680 ;
    END
  END gpio_in[4]
  PIN gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 559.000 2600.000 559.600 ;
    END
  END gpio_in[5]
  PIN gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 656.920 2600.000 657.520 ;
    END
  END gpio_in[6]
  PIN gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 754.840 2600.000 755.440 ;
    END
  END gpio_in[7]
  PIN gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 852.760 2600.000 853.360 ;
    END
  END gpio_in[8]
  PIN gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 950.680 2600.000 951.280 ;
    END
  END gpio_in[9]
  PIN gpio_loopback_one[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2597.600 151.000 2600.000 151.600 ;
    END
  END gpio_loopback_one[0]
  PIN gpio_loopback_one[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1130.200 2600.000 1130.800 ;
    END
  END gpio_loopback_one[10]
  PIN gpio_loopback_one[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1228.120 2600.000 1228.720 ;
    END
  END gpio_loopback_one[11]
  PIN gpio_loopback_one[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1326.040 2600.000 1326.640 ;
    END
  END gpio_loopback_one[12]
  PIN gpio_loopback_one[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1423.960 2600.000 1424.560 ;
    END
  END gpio_loopback_one[13]
  PIN gpio_loopback_one[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1521.880 2600.000 1522.480 ;
    END
  END gpio_loopback_one[14]
  PIN gpio_loopback_one[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2340.110 1597.600 2340.390 1600.000 ;
    END
  END gpio_loopback_one[15]
  PIN gpio_loopback_one[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.070 1597.600 2053.350 1600.000 ;
    END
  END gpio_loopback_one[16]
  PIN gpio_loopback_one[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 1597.600 1766.310 1600.000 ;
    END
  END gpio_loopback_one[17]
  PIN gpio_loopback_one[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 1597.600 1479.270 1600.000 ;
    END
  END gpio_loopback_one[18]
  PIN gpio_loopback_one[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 1597.600 1192.230 1600.000 ;
    END
  END gpio_loopback_one[19]
  PIN gpio_loopback_one[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 248.920 2600.000 249.520 ;
    END
  END gpio_loopback_one[1]
  PIN gpio_loopback_one[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 1597.600 905.190 1600.000 ;
    END
  END gpio_loopback_one[20]
  PIN gpio_loopback_one[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 1597.600 618.150 1600.000 ;
    END
  END gpio_loopback_one[21]
  PIN gpio_loopback_one[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 1597.600 331.110 1600.000 ;
    END
  END gpio_loopback_one[22]
  PIN gpio_loopback_one[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 1597.600 44.070 1600.000 ;
    END
  END gpio_loopback_one[23]
  PIN gpio_loopback_one[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 2.400 1408.240 ;
    END
  END gpio_loopback_one[24]
  PIN gpio_loopback_one[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.720 2.400 1310.320 ;
    END
  END gpio_loopback_one[25]
  PIN gpio_loopback_one[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1211.800 2.400 1212.400 ;
    END
  END gpio_loopback_one[26]
  PIN gpio_loopback_one[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.880 2.400 1114.480 ;
    END
  END gpio_loopback_one[27]
  PIN gpio_loopback_one[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.960 2.400 1016.560 ;
    END
  END gpio_loopback_one[28]
  PIN gpio_loopback_one[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 2.400 918.640 ;
    END
  END gpio_loopback_one[29]
  PIN gpio_loopback_one[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 346.840 2600.000 347.440 ;
    END
  END gpio_loopback_one[2]
  PIN gpio_loopback_one[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 2.400 820.720 ;
    END
  END gpio_loopback_one[30]
  PIN gpio_loopback_one[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 2.400 722.800 ;
    END
  END gpio_loopback_one[31]
  PIN gpio_loopback_one[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 2.400 624.880 ;
    END
  END gpio_loopback_one[32]
  PIN gpio_loopback_one[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 2.400 526.960 ;
    END
  END gpio_loopback_one[33]
  PIN gpio_loopback_one[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 2.400 429.040 ;
    END
  END gpio_loopback_one[34]
  PIN gpio_loopback_one[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 2.400 331.120 ;
    END
  END gpio_loopback_one[35]
  PIN gpio_loopback_one[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 2.400 233.200 ;
    END
  END gpio_loopback_one[36]
  PIN gpio_loopback_one[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 2.400 135.280 ;
    END
  END gpio_loopback_one[37]
  PIN gpio_loopback_one[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 2.400 ;
    END
  END gpio_loopback_one[38]
  PIN gpio_loopback_one[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 2.400 ;
    END
  END gpio_loopback_one[39]
  PIN gpio_loopback_one[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 444.760 2600.000 445.360 ;
    END
  END gpio_loopback_one[3]
  PIN gpio_loopback_one[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 2.400 ;
    END
  END gpio_loopback_one[40]
  PIN gpio_loopback_one[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 0.000 1177.970 2.400 ;
    END
  END gpio_loopback_one[41]
  PIN gpio_loopback_one[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.250 0.000 1470.530 2.400 ;
    END
  END gpio_loopback_one[42]
  PIN gpio_loopback_one[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.810 0.000 1763.090 2.400 ;
    END
  END gpio_loopback_one[43]
  PIN gpio_loopback_one[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 542.680 2600.000 543.280 ;
    END
  END gpio_loopback_one[4]
  PIN gpio_loopback_one[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 640.600 2600.000 641.200 ;
    END
  END gpio_loopback_one[5]
  PIN gpio_loopback_one[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 738.520 2600.000 739.120 ;
    END
  END gpio_loopback_one[6]
  PIN gpio_loopback_one[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 836.440 2600.000 837.040 ;
    END
  END gpio_loopback_one[7]
  PIN gpio_loopback_one[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 934.360 2600.000 934.960 ;
    END
  END gpio_loopback_one[8]
  PIN gpio_loopback_one[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1032.280 2600.000 1032.880 ;
    END
  END gpio_loopback_one[9]
  PIN gpio_loopback_zero[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2597.600 159.160 2600.000 159.760 ;
    END
  END gpio_loopback_zero[0]
  PIN gpio_loopback_zero[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1138.360 2600.000 1138.960 ;
    END
  END gpio_loopback_zero[10]
  PIN gpio_loopback_zero[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1236.280 2600.000 1236.880 ;
    END
  END gpio_loopback_zero[11]
  PIN gpio_loopback_zero[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1334.200 2600.000 1334.800 ;
    END
  END gpio_loopback_zero[12]
  PIN gpio_loopback_zero[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1432.120 2600.000 1432.720 ;
    END
  END gpio_loopback_zero[13]
  PIN gpio_loopback_zero[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1530.040 2600.000 1530.640 ;
    END
  END gpio_loopback_zero[14]
  PIN gpio_loopback_zero[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 2316.190 1597.600 2316.470 1600.000 ;
    END
  END gpio_loopback_zero[15]
  PIN gpio_loopback_zero[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.150 1597.600 2029.430 1600.000 ;
    END
  END gpio_loopback_zero[16]
  PIN gpio_loopback_zero[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.110 1597.600 1742.390 1600.000 ;
    END
  END gpio_loopback_zero[17]
  PIN gpio_loopback_zero[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 1597.600 1455.350 1600.000 ;
    END
  END gpio_loopback_zero[18]
  PIN gpio_loopback_zero[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 1597.600 1168.310 1600.000 ;
    END
  END gpio_loopback_zero[19]
  PIN gpio_loopback_zero[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2597.600 257.080 2600.000 257.680 ;
    END
  END gpio_loopback_zero[1]
  PIN gpio_loopback_zero[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 1597.600 881.270 1600.000 ;
    END
  END gpio_loopback_zero[20]
  PIN gpio_loopback_zero[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1597.600 594.230 1600.000 ;
    END
  END gpio_loopback_zero[21]
  PIN gpio_loopback_zero[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 1597.600 307.190 1600.000 ;
    END
  END gpio_loopback_zero[22]
  PIN gpio_loopback_zero[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 1597.600 20.150 1600.000 ;
    END
  END gpio_loopback_zero[23]
  PIN gpio_loopback_zero[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1399.480 2.400 1400.080 ;
    END
  END gpio_loopback_zero[24]
  PIN gpio_loopback_zero[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1301.560 2.400 1302.160 ;
    END
  END gpio_loopback_zero[25]
  PIN gpio_loopback_zero[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1203.640 2.400 1204.240 ;
    END
  END gpio_loopback_zero[26]
  PIN gpio_loopback_zero[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.720 2.400 1106.320 ;
    END
  END gpio_loopback_zero[27]
  PIN gpio_loopback_zero[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 2.400 1008.400 ;
    END
  END gpio_loopback_zero[28]
  PIN gpio_loopback_zero[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 2.400 910.480 ;
    END
  END gpio_loopback_zero[29]
  PIN gpio_loopback_zero[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 355.000 2600.000 355.600 ;
    END
  END gpio_loopback_zero[2]
  PIN gpio_loopback_zero[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 2.400 812.560 ;
    END
  END gpio_loopback_zero[30]
  PIN gpio_loopback_zero[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 2.400 714.640 ;
    END
  END gpio_loopback_zero[31]
  PIN gpio_loopback_zero[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 2.400 616.720 ;
    END
  END gpio_loopback_zero[32]
  PIN gpio_loopback_zero[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 2.400 518.800 ;
    END
  END gpio_loopback_zero[33]
  PIN gpio_loopback_zero[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 2.400 420.880 ;
    END
  END gpio_loopback_zero[34]
  PIN gpio_loopback_zero[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 2.400 322.960 ;
    END
  END gpio_loopback_zero[35]
  PIN gpio_loopback_zero[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 2.400 225.040 ;
    END
  END gpio_loopback_zero[36]
  PIN gpio_loopback_zero[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END gpio_loopback_zero[37]
  PIN gpio_loopback_zero[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 2.400 ;
    END
  END gpio_loopback_zero[38]
  PIN gpio_loopback_zero[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 2.400 ;
    END
  END gpio_loopback_zero[39]
  PIN gpio_loopback_zero[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 452.920 2600.000 453.520 ;
    END
  END gpio_loopback_zero[3]
  PIN gpio_loopback_zero[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 2.400 ;
    END
  END gpio_loopback_zero[40]
  PIN gpio_loopback_zero[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 0.000 1202.350 2.400 ;
    END
  END gpio_loopback_zero[41]
  PIN gpio_loopback_zero[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.630 0.000 1494.910 2.400 ;
    END
  END gpio_loopback_zero[42]
  PIN gpio_loopback_zero[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 2.400 ;
    END
  END gpio_loopback_zero[43]
  PIN gpio_loopback_zero[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 550.840 2600.000 551.440 ;
    END
  END gpio_loopback_zero[4]
  PIN gpio_loopback_zero[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 648.760 2600.000 649.360 ;
    END
  END gpio_loopback_zero[5]
  PIN gpio_loopback_zero[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 746.680 2600.000 747.280 ;
    END
  END gpio_loopback_zero[6]
  PIN gpio_loopback_zero[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 844.600 2600.000 845.200 ;
    END
  END gpio_loopback_zero[7]
  PIN gpio_loopback_zero[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 942.520 2600.000 943.120 ;
    END
  END gpio_loopback_zero[8]
  PIN gpio_loopback_zero[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1040.440 2600.000 1041.040 ;
    END
  END gpio_loopback_zero[9]
  PIN gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 142.840 2600.000 143.440 ;
    END
  END gpio_oeb[0]
  PIN gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1122.040 2600.000 1122.640 ;
    END
  END gpio_oeb[10]
  PIN gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1219.960 2600.000 1220.560 ;
    END
  END gpio_oeb[11]
  PIN gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1317.880 2600.000 1318.480 ;
    END
  END gpio_oeb[12]
  PIN gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1415.800 2600.000 1416.400 ;
    END
  END gpio_oeb[13]
  PIN gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1513.720 2600.000 1514.320 ;
    END
  END gpio_oeb[14]
  PIN gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2364.030 1597.600 2364.310 1600.000 ;
    END
  END gpio_oeb[15]
  PIN gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2076.990 1597.600 2077.270 1600.000 ;
    END
  END gpio_oeb[16]
  PIN gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1789.950 1597.600 1790.230 1600.000 ;
    END
  END gpio_oeb[17]
  PIN gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1502.910 1597.600 1503.190 1600.000 ;
    END
  END gpio_oeb[18]
  PIN gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1215.870 1597.600 1216.150 1600.000 ;
    END
  END gpio_oeb[19]
  PIN gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 240.760 2600.000 241.360 ;
    END
  END gpio_oeb[1]
  PIN gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 928.830 1597.600 929.110 1600.000 ;
    END
  END gpio_oeb[20]
  PIN gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 641.790 1597.600 642.070 1600.000 ;
    END
  END gpio_oeb[21]
  PIN gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 354.750 1597.600 355.030 1600.000 ;
    END
  END gpio_oeb[22]
  PIN gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 67.710 1597.600 67.990 1600.000 ;
    END
  END gpio_oeb[23]
  PIN gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1415.800 2.400 1416.400 ;
    END
  END gpio_oeb[24]
  PIN gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.880 2.400 1318.480 ;
    END
  END gpio_oeb[25]
  PIN gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1219.960 2.400 1220.560 ;
    END
  END gpio_oeb[26]
  PIN gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 2.400 1122.640 ;
    END
  END gpio_oeb[27]
  PIN gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 2.400 1024.720 ;
    END
  END gpio_oeb[28]
  PIN gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 2.400 926.800 ;
    END
  END gpio_oeb[29]
  PIN gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 338.680 2600.000 339.280 ;
    END
  END gpio_oeb[2]
  PIN gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 2.400 828.880 ;
    END
  END gpio_oeb[30]
  PIN gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 2.400 730.960 ;
    END
  END gpio_oeb[31]
  PIN gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 2.400 633.040 ;
    END
  END gpio_oeb[32]
  PIN gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 2.400 535.120 ;
    END
  END gpio_oeb[33]
  PIN gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 2.400 437.200 ;
    END
  END gpio_oeb[34]
  PIN gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 2.400 339.280 ;
    END
  END gpio_oeb[35]
  PIN gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 2.400 241.360 ;
    END
  END gpio_oeb[36]
  PIN gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 2.400 143.440 ;
    END
  END gpio_oeb[37]
  PIN gpio_oeb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 2.400 ;
    END
  END gpio_oeb[38]
  PIN gpio_oeb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 2.400 ;
    END
  END gpio_oeb[39]
  PIN gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 436.600 2600.000 437.200 ;
    END
  END gpio_oeb[3]
  PIN gpio_oeb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 2.400 ;
    END
  END gpio_oeb[40]
  PIN gpio_oeb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 2.400 ;
    END
  END gpio_oeb[41]
  PIN gpio_oeb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 2.400 ;
    END
  END gpio_oeb[42]
  PIN gpio_oeb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1738.430 0.000 1738.710 2.400 ;
    END
  END gpio_oeb[43]
  PIN gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 534.520 2600.000 535.120 ;
    END
  END gpio_oeb[4]
  PIN gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 632.440 2600.000 633.040 ;
    END
  END gpio_oeb[5]
  PIN gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 730.360 2600.000 730.960 ;
    END
  END gpio_oeb[6]
  PIN gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 828.280 2600.000 828.880 ;
    END
  END gpio_oeb[7]
  PIN gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 926.200 2600.000 926.800 ;
    END
  END gpio_oeb[8]
  PIN gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1024.120 2600.000 1024.720 ;
    END
  END gpio_oeb[9]
  PIN gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 118.360 2600.000 118.960 ;
    END
  END gpio_out[0]
  PIN gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1097.560 2600.000 1098.160 ;
    END
  END gpio_out[10]
  PIN gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1195.480 2600.000 1196.080 ;
    END
  END gpio_out[11]
  PIN gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1293.400 2600.000 1294.000 ;
    END
  END gpio_out[12]
  PIN gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1391.320 2600.000 1391.920 ;
    END
  END gpio_out[13]
  PIN gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1489.240 2600.000 1489.840 ;
    END
  END gpio_out[14]
  PIN gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2435.790 1597.600 2436.070 1600.000 ;
    END
  END gpio_out[15]
  PIN gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2148.750 1597.600 2149.030 1600.000 ;
    END
  END gpio_out[16]
  PIN gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1861.710 1597.600 1861.990 1600.000 ;
    END
  END gpio_out[17]
  PIN gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1574.670 1597.600 1574.950 1600.000 ;
    END
  END gpio_out[18]
  PIN gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1287.630 1597.600 1287.910 1600.000 ;
    END
  END gpio_out[19]
  PIN gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 216.280 2600.000 216.880 ;
    END
  END gpio_out[1]
  PIN gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1000.590 1597.600 1000.870 1600.000 ;
    END
  END gpio_out[20]
  PIN gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 713.550 1597.600 713.830 1600.000 ;
    END
  END gpio_out[21]
  PIN gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 426.510 1597.600 426.790 1600.000 ;
    END
  END gpio_out[22]
  PIN gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 139.470 1597.600 139.750 1600.000 ;
    END
  END gpio_out[23]
  PIN gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.280 2.400 1440.880 ;
    END
  END gpio_out[24]
  PIN gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 2.400 1342.960 ;
    END
  END gpio_out[25]
  PIN gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 2.400 1245.040 ;
    END
  END gpio_out[26]
  PIN gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1146.520 2.400 1147.120 ;
    END
  END gpio_out[27]
  PIN gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 2.400 1049.200 ;
    END
  END gpio_out[28]
  PIN gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 2.400 951.280 ;
    END
  END gpio_out[29]
  PIN gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 314.200 2600.000 314.800 ;
    END
  END gpio_out[2]
  PIN gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.760 2.400 853.360 ;
    END
  END gpio_out[30]
  PIN gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 2.400 755.440 ;
    END
  END gpio_out[31]
  PIN gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 2.400 657.520 ;
    END
  END gpio_out[32]
  PIN gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 2.400 559.600 ;
    END
  END gpio_out[33]
  PIN gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 2.400 461.680 ;
    END
  END gpio_out[34]
  PIN gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 2.400 363.760 ;
    END
  END gpio_out[35]
  PIN gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 2.400 265.840 ;
    END
  END gpio_out[36]
  PIN gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 2.400 167.920 ;
    END
  END gpio_out[37]
  PIN gpio_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 2.400 ;
    END
  END gpio_out[38]
  PIN gpio_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 2.400 ;
    END
  END gpio_out[39]
  PIN gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 412.120 2600.000 412.720 ;
    END
  END gpio_out[3]
  PIN gpio_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.397600 ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 2.400 ;
    END
  END gpio_out[40]
  PIN gpio_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 2.400 ;
    END
  END gpio_out[41]
  PIN gpio_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 2.400 ;
    END
  END gpio_out[42]
  PIN gpio_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1665.290 0.000 1665.570 2.400 ;
    END
  END gpio_out[43]
  PIN gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 510.040 2600.000 510.640 ;
    END
  END gpio_out[4]
  PIN gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 607.960 2600.000 608.560 ;
    END
  END gpio_out[5]
  PIN gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 705.880 2600.000 706.480 ;
    END
  END gpio_out[6]
  PIN gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 803.800 2600.000 804.400 ;
    END
  END gpio_out[7]
  PIN gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 901.720 2600.000 902.320 ;
    END
  END gpio_out[8]
  PIN gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 999.640 2600.000 1000.240 ;
    END
  END gpio_out[9]
  PIN gpio_slow_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 77.560 2600.000 78.160 ;
    END
  END gpio_slow_sel[0]
  PIN gpio_slow_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1056.760 2600.000 1057.360 ;
    END
  END gpio_slow_sel[10]
  PIN gpio_slow_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1154.680 2600.000 1155.280 ;
    END
  END gpio_slow_sel[11]
  PIN gpio_slow_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1252.600 2600.000 1253.200 ;
    END
  END gpio_slow_sel[12]
  PIN gpio_slow_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1350.520 2600.000 1351.120 ;
    END
  END gpio_slow_sel[13]
  PIN gpio_slow_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1448.440 2600.000 1449.040 ;
    END
  END gpio_slow_sel[14]
  PIN gpio_slow_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2555.390 1597.600 2555.670 1600.000 ;
    END
  END gpio_slow_sel[15]
  PIN gpio_slow_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2268.350 1597.600 2268.630 1600.000 ;
    END
  END gpio_slow_sel[16]
  PIN gpio_slow_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1981.310 1597.600 1981.590 1600.000 ;
    END
  END gpio_slow_sel[17]
  PIN gpio_slow_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1694.270 1597.600 1694.550 1600.000 ;
    END
  END gpio_slow_sel[18]
  PIN gpio_slow_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1407.230 1597.600 1407.510 1600.000 ;
    END
  END gpio_slow_sel[19]
  PIN gpio_slow_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 175.480 2600.000 176.080 ;
    END
  END gpio_slow_sel[1]
  PIN gpio_slow_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1120.190 1597.600 1120.470 1600.000 ;
    END
  END gpio_slow_sel[20]
  PIN gpio_slow_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 833.150 1597.600 833.430 1600.000 ;
    END
  END gpio_slow_sel[21]
  PIN gpio_slow_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 546.110 1597.600 546.390 1600.000 ;
    END
  END gpio_slow_sel[22]
  PIN gpio_slow_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 259.070 1597.600 259.350 1600.000 ;
    END
  END gpio_slow_sel[23]
  PIN gpio_slow_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1481.080 2.400 1481.680 ;
    END
  END gpio_slow_sel[24]
  PIN gpio_slow_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.160 2.400 1383.760 ;
    END
  END gpio_slow_sel[25]
  PIN gpio_slow_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 2.400 1285.840 ;
    END
  END gpio_slow_sel[26]
  PIN gpio_slow_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1187.320 2.400 1187.920 ;
    END
  END gpio_slow_sel[27]
  PIN gpio_slow_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1089.400 2.400 1090.000 ;
    END
  END gpio_slow_sel[28]
  PIN gpio_slow_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 2.400 992.080 ;
    END
  END gpio_slow_sel[29]
  PIN gpio_slow_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 273.400 2600.000 274.000 ;
    END
  END gpio_slow_sel[2]
  PIN gpio_slow_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 2.400 894.160 ;
    END
  END gpio_slow_sel[30]
  PIN gpio_slow_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 2.400 796.240 ;
    END
  END gpio_slow_sel[31]
  PIN gpio_slow_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 2.400 698.320 ;
    END
  END gpio_slow_sel[32]
  PIN gpio_slow_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 2.400 600.400 ;
    END
  END gpio_slow_sel[33]
  PIN gpio_slow_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 2.400 502.480 ;
    END
  END gpio_slow_sel[34]
  PIN gpio_slow_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 2.400 404.560 ;
    END
  END gpio_slow_sel[35]
  PIN gpio_slow_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 2.400 306.640 ;
    END
  END gpio_slow_sel[36]
  PIN gpio_slow_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 2.400 208.720 ;
    END
  END gpio_slow_sel[37]
  PIN gpio_slow_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END gpio_slow_sel[38]
  PIN gpio_slow_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 2.400 ;
    END
  END gpio_slow_sel[39]
  PIN gpio_slow_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 371.320 2600.000 371.920 ;
    END
  END gpio_slow_sel[3]
  PIN gpio_slow_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 2.400 ;
    END
  END gpio_slow_sel[40]
  PIN gpio_slow_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 2.400 ;
    END
  END gpio_slow_sel[41]
  PIN gpio_slow_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1250.830 0.000 1251.110 2.400 ;
    END
  END gpio_slow_sel[42]
  PIN gpio_slow_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1543.390 0.000 1543.670 2.400 ;
    END
  END gpio_slow_sel[43]
  PIN gpio_slow_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 469.240 2600.000 469.840 ;
    END
  END gpio_slow_sel[4]
  PIN gpio_slow_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 567.160 2600.000 567.760 ;
    END
  END gpio_slow_sel[5]
  PIN gpio_slow_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 665.080 2600.000 665.680 ;
    END
  END gpio_slow_sel[6]
  PIN gpio_slow_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 763.000 2600.000 763.600 ;
    END
  END gpio_slow_sel[7]
  PIN gpio_slow_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 860.920 2600.000 861.520 ;
    END
  END gpio_slow_sel[8]
  PIN gpio_slow_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 958.840 2600.000 959.440 ;
    END
  END gpio_slow_sel[9]
  PIN gpio_vtrip_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 126.520 2600.000 127.120 ;
    END
  END gpio_vtrip_sel[0]
  PIN gpio_vtrip_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1105.720 2600.000 1106.320 ;
    END
  END gpio_vtrip_sel[10]
  PIN gpio_vtrip_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1203.640 2600.000 1204.240 ;
    END
  END gpio_vtrip_sel[11]
  PIN gpio_vtrip_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1301.560 2600.000 1302.160 ;
    END
  END gpio_vtrip_sel[12]
  PIN gpio_vtrip_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1399.480 2600.000 1400.080 ;
    END
  END gpio_vtrip_sel[13]
  PIN gpio_vtrip_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1497.400 2600.000 1498.000 ;
    END
  END gpio_vtrip_sel[14]
  PIN gpio_vtrip_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2411.870 1597.600 2412.150 1600.000 ;
    END
  END gpio_vtrip_sel[15]
  PIN gpio_vtrip_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 2124.830 1597.600 2125.110 1600.000 ;
    END
  END gpio_vtrip_sel[16]
  PIN gpio_vtrip_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1837.790 1597.600 1838.070 1600.000 ;
    END
  END gpio_vtrip_sel[17]
  PIN gpio_vtrip_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1550.750 1597.600 1551.030 1600.000 ;
    END
  END gpio_vtrip_sel[18]
  PIN gpio_vtrip_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1263.710 1597.600 1263.990 1600.000 ;
    END
  END gpio_vtrip_sel[19]
  PIN gpio_vtrip_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 224.440 2600.000 225.040 ;
    END
  END gpio_vtrip_sel[1]
  PIN gpio_vtrip_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 976.670 1597.600 976.950 1600.000 ;
    END
  END gpio_vtrip_sel[20]
  PIN gpio_vtrip_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 689.630 1597.600 689.910 1600.000 ;
    END
  END gpio_vtrip_sel[21]
  PIN gpio_vtrip_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 402.590 1597.600 402.870 1600.000 ;
    END
  END gpio_vtrip_sel[22]
  PIN gpio_vtrip_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 115.550 1597.600 115.830 1600.000 ;
    END
  END gpio_vtrip_sel[23]
  PIN gpio_vtrip_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1432.120 2.400 1432.720 ;
    END
  END gpio_vtrip_sel[24]
  PIN gpio_vtrip_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1334.200 2.400 1334.800 ;
    END
  END gpio_vtrip_sel[25]
  PIN gpio_vtrip_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 2.400 1236.880 ;
    END
  END gpio_vtrip_sel[26]
  PIN gpio_vtrip_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1138.360 2.400 1138.960 ;
    END
  END gpio_vtrip_sel[27]
  PIN gpio_vtrip_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 2.400 1041.040 ;
    END
  END gpio_vtrip_sel[28]
  PIN gpio_vtrip_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 942.520 2.400 943.120 ;
    END
  END gpio_vtrip_sel[29]
  PIN gpio_vtrip_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 322.360 2600.000 322.960 ;
    END
  END gpio_vtrip_sel[2]
  PIN gpio_vtrip_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 2.400 845.200 ;
    END
  END gpio_vtrip_sel[30]
  PIN gpio_vtrip_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 2.400 747.280 ;
    END
  END gpio_vtrip_sel[31]
  PIN gpio_vtrip_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 2.400 649.360 ;
    END
  END gpio_vtrip_sel[32]
  PIN gpio_vtrip_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 2.400 551.440 ;
    END
  END gpio_vtrip_sel[33]
  PIN gpio_vtrip_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 2.400 453.520 ;
    END
  END gpio_vtrip_sel[34]
  PIN gpio_vtrip_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 2.400 355.600 ;
    END
  END gpio_vtrip_sel[35]
  PIN gpio_vtrip_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 2.400 257.680 ;
    END
  END gpio_vtrip_sel[36]
  PIN gpio_vtrip_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 2.400 159.760 ;
    END
  END gpio_vtrip_sel[37]
  PIN gpio_vtrip_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 2.400 ;
    END
  END gpio_vtrip_sel[38]
  PIN gpio_vtrip_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 2.400 ;
    END
  END gpio_vtrip_sel[39]
  PIN gpio_vtrip_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 420.280 2600.000 420.880 ;
    END
  END gpio_vtrip_sel[3]
  PIN gpio_vtrip_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 2.400 ;
    END
  END gpio_vtrip_sel[40]
  PIN gpio_vtrip_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 2.400 ;
    END
  END gpio_vtrip_sel[41]
  PIN gpio_vtrip_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 2.400 ;
    END
  END gpio_vtrip_sel[42]
  PIN gpio_vtrip_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 1689.670 0.000 1689.950 2.400 ;
    END
  END gpio_vtrip_sel[43]
  PIN gpio_vtrip_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 518.200 2600.000 518.800 ;
    END
  END gpio_vtrip_sel[4]
  PIN gpio_vtrip_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 616.120 2600.000 616.720 ;
    END
  END gpio_vtrip_sel[5]
  PIN gpio_vtrip_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 714.040 2600.000 714.640 ;
    END
  END gpio_vtrip_sel[6]
  PIN gpio_vtrip_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 811.960 2600.000 812.560 ;
    END
  END gpio_vtrip_sel[7]
  PIN gpio_vtrip_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 909.880 2600.000 910.480 ;
    END
  END gpio_vtrip_sel[8]
  PIN gpio_vtrip_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 2597.600 1007.800 2600.000 1008.400 ;
    END
  END gpio_vtrip_sel[9]
  PIN mask_rev[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1811.570 0.000 1811.850 2.400 ;
    END
  END mask_rev[0]
  PIN mask_rev[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2055.370 0.000 2055.650 2.400 ;
    END
  END mask_rev[10]
  PIN mask_rev[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2079.750 0.000 2080.030 2.400 ;
    END
  END mask_rev[11]
  PIN mask_rev[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2104.130 0.000 2104.410 2.400 ;
    END
  END mask_rev[12]
  PIN mask_rev[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2128.510 0.000 2128.790 2.400 ;
    END
  END mask_rev[13]
  PIN mask_rev[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2152.890 0.000 2153.170 2.400 ;
    END
  END mask_rev[14]
  PIN mask_rev[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2177.270 0.000 2177.550 2.400 ;
    END
  END mask_rev[15]
  PIN mask_rev[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2201.650 0.000 2201.930 2.400 ;
    END
  END mask_rev[16]
  PIN mask_rev[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2226.030 0.000 2226.310 2.400 ;
    END
  END mask_rev[17]
  PIN mask_rev[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 2250.410 0.000 2250.690 2.400 ;
    END
  END mask_rev[18]
  PIN mask_rev[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2274.790 0.000 2275.070 2.400 ;
    END
  END mask_rev[19]
  PIN mask_rev[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1835.950 0.000 1836.230 2.400 ;
    END
  END mask_rev[1]
  PIN mask_rev[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 2299.170 0.000 2299.450 2.400 ;
    END
  END mask_rev[20]
  PIN mask_rev[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 2323.550 0.000 2323.830 2.400 ;
    END
  END mask_rev[21]
  PIN mask_rev[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 2347.930 0.000 2348.210 2.400 ;
    END
  END mask_rev[22]
  PIN mask_rev[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 2372.310 0.000 2372.590 2.400 ;
    END
  END mask_rev[23]
  PIN mask_rev[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2396.690 0.000 2396.970 2.400 ;
    END
  END mask_rev[24]
  PIN mask_rev[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2421.070 0.000 2421.350 2.400 ;
    END
  END mask_rev[25]
  PIN mask_rev[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2445.450 0.000 2445.730 2.400 ;
    END
  END mask_rev[26]
  PIN mask_rev[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2469.830 0.000 2470.110 2.400 ;
    END
  END mask_rev[27]
  PIN mask_rev[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2494.210 0.000 2494.490 2.400 ;
    END
  END mask_rev[28]
  PIN mask_rev[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2518.590 0.000 2518.870 2.400 ;
    END
  END mask_rev[29]
  PIN mask_rev[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1860.330 0.000 1860.610 2.400 ;
    END
  END mask_rev[2]
  PIN mask_rev[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2542.970 0.000 2543.250 2.400 ;
    END
  END mask_rev[30]
  PIN mask_rev[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2567.350 0.000 2567.630 2.400 ;
    END
  END mask_rev[31]
  PIN mask_rev[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1884.710 0.000 1884.990 2.400 ;
    END
  END mask_rev[3]
  PIN mask_rev[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1909.090 0.000 1909.370 2.400 ;
    END
  END mask_rev[4]
  PIN mask_rev[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1933.470 0.000 1933.750 2.400 ;
    END
  END mask_rev[5]
  PIN mask_rev[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 1957.850 0.000 1958.130 2.400 ;
    END
  END mask_rev[6]
  PIN mask_rev[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1982.230 0.000 1982.510 2.400 ;
    END
  END mask_rev[7]
  PIN mask_rev[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2006.610 0.000 2006.890 2.400 ;
    END
  END mask_rev[8]
  PIN mask_rev[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2030.990 0.000 2031.270 2.400 ;
    END
  END mask_rev[9]
  PIN por
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END por
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END porb
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END resetb
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2594.400 1588.565 ;
      LAYER met1 ;
        RECT 0.070 9.560 2599.850 1591.840 ;
      LAYER met2 ;
        RECT 0.090 1597.320 19.590 1598.410 ;
        RECT 20.430 1597.320 43.510 1598.410 ;
        RECT 44.350 1597.320 67.430 1598.410 ;
        RECT 68.270 1597.320 91.350 1598.410 ;
        RECT 92.190 1597.320 115.270 1598.410 ;
        RECT 116.110 1597.320 139.190 1598.410 ;
        RECT 140.030 1597.320 163.110 1598.410 ;
        RECT 163.950 1597.320 187.030 1598.410 ;
        RECT 187.870 1597.320 210.950 1598.410 ;
        RECT 211.790 1597.320 234.870 1598.410 ;
        RECT 235.710 1597.320 258.790 1598.410 ;
        RECT 259.630 1597.320 282.710 1598.410 ;
        RECT 283.550 1597.320 306.630 1598.410 ;
        RECT 307.470 1597.320 330.550 1598.410 ;
        RECT 331.390 1597.320 354.470 1598.410 ;
        RECT 355.310 1597.320 378.390 1598.410 ;
        RECT 379.230 1597.320 402.310 1598.410 ;
        RECT 403.150 1597.320 426.230 1598.410 ;
        RECT 427.070 1597.320 450.150 1598.410 ;
        RECT 450.990 1597.320 474.070 1598.410 ;
        RECT 474.910 1597.320 497.990 1598.410 ;
        RECT 498.830 1597.320 521.910 1598.410 ;
        RECT 522.750 1597.320 545.830 1598.410 ;
        RECT 546.670 1597.320 569.750 1598.410 ;
        RECT 570.590 1597.320 593.670 1598.410 ;
        RECT 594.510 1597.320 617.590 1598.410 ;
        RECT 618.430 1597.320 641.510 1598.410 ;
        RECT 642.350 1597.320 665.430 1598.410 ;
        RECT 666.270 1597.320 689.350 1598.410 ;
        RECT 690.190 1597.320 713.270 1598.410 ;
        RECT 714.110 1597.320 737.190 1598.410 ;
        RECT 738.030 1597.320 761.110 1598.410 ;
        RECT 761.950 1597.320 785.030 1598.410 ;
        RECT 785.870 1597.320 808.950 1598.410 ;
        RECT 809.790 1597.320 832.870 1598.410 ;
        RECT 833.710 1597.320 856.790 1598.410 ;
        RECT 857.630 1597.320 880.710 1598.410 ;
        RECT 881.550 1597.320 904.630 1598.410 ;
        RECT 905.470 1597.320 928.550 1598.410 ;
        RECT 929.390 1597.320 952.470 1598.410 ;
        RECT 953.310 1597.320 976.390 1598.410 ;
        RECT 977.230 1597.320 1000.310 1598.410 ;
        RECT 1001.150 1597.320 1024.230 1598.410 ;
        RECT 1025.070 1597.320 1048.150 1598.410 ;
        RECT 1048.990 1597.320 1072.070 1598.410 ;
        RECT 1072.910 1597.320 1095.990 1598.410 ;
        RECT 1096.830 1597.320 1119.910 1598.410 ;
        RECT 1120.750 1597.320 1143.830 1598.410 ;
        RECT 1144.670 1597.320 1167.750 1598.410 ;
        RECT 1168.590 1597.320 1191.670 1598.410 ;
        RECT 1192.510 1597.320 1215.590 1598.410 ;
        RECT 1216.430 1597.320 1239.510 1598.410 ;
        RECT 1240.350 1597.320 1263.430 1598.410 ;
        RECT 1264.270 1597.320 1287.350 1598.410 ;
        RECT 1288.190 1597.320 1311.270 1598.410 ;
        RECT 1312.110 1597.320 1335.190 1598.410 ;
        RECT 1336.030 1597.320 1359.110 1598.410 ;
        RECT 1359.950 1597.320 1383.030 1598.410 ;
        RECT 1383.870 1597.320 1406.950 1598.410 ;
        RECT 1407.790 1597.320 1430.870 1598.410 ;
        RECT 1431.710 1597.320 1454.790 1598.410 ;
        RECT 1455.630 1597.320 1478.710 1598.410 ;
        RECT 1479.550 1597.320 1502.630 1598.410 ;
        RECT 1503.470 1597.320 1526.550 1598.410 ;
        RECT 1527.390 1597.320 1550.470 1598.410 ;
        RECT 1551.310 1597.320 1574.390 1598.410 ;
        RECT 1575.230 1597.320 1598.310 1598.410 ;
        RECT 1599.150 1597.320 1622.230 1598.410 ;
        RECT 1623.070 1597.320 1646.150 1598.410 ;
        RECT 1646.990 1597.320 1670.070 1598.410 ;
        RECT 1670.910 1597.320 1693.990 1598.410 ;
        RECT 1694.830 1597.320 1717.910 1598.410 ;
        RECT 1718.750 1597.320 1741.830 1598.410 ;
        RECT 1742.670 1597.320 1765.750 1598.410 ;
        RECT 1766.590 1597.320 1789.670 1598.410 ;
        RECT 1790.510 1597.320 1813.590 1598.410 ;
        RECT 1814.430 1597.320 1837.510 1598.410 ;
        RECT 1838.350 1597.320 1861.430 1598.410 ;
        RECT 1862.270 1597.320 1885.350 1598.410 ;
        RECT 1886.190 1597.320 1909.270 1598.410 ;
        RECT 1910.110 1597.320 1933.190 1598.410 ;
        RECT 1934.030 1597.320 1957.110 1598.410 ;
        RECT 1957.950 1597.320 1981.030 1598.410 ;
        RECT 1981.870 1597.320 2004.950 1598.410 ;
        RECT 2005.790 1597.320 2028.870 1598.410 ;
        RECT 2029.710 1597.320 2052.790 1598.410 ;
        RECT 2053.630 1597.320 2076.710 1598.410 ;
        RECT 2077.550 1597.320 2100.630 1598.410 ;
        RECT 2101.470 1597.320 2124.550 1598.410 ;
        RECT 2125.390 1597.320 2148.470 1598.410 ;
        RECT 2149.310 1597.320 2172.390 1598.410 ;
        RECT 2173.230 1597.320 2196.310 1598.410 ;
        RECT 2197.150 1597.320 2220.230 1598.410 ;
        RECT 2221.070 1597.320 2244.150 1598.410 ;
        RECT 2244.990 1597.320 2268.070 1598.410 ;
        RECT 2268.910 1597.320 2291.990 1598.410 ;
        RECT 2292.830 1597.320 2315.910 1598.410 ;
        RECT 2316.750 1597.320 2339.830 1598.410 ;
        RECT 2340.670 1597.320 2363.750 1598.410 ;
        RECT 2364.590 1597.320 2387.670 1598.410 ;
        RECT 2388.510 1597.320 2411.590 1598.410 ;
        RECT 2412.430 1597.320 2435.510 1598.410 ;
        RECT 2436.350 1597.320 2459.430 1598.410 ;
        RECT 2460.270 1597.320 2483.350 1598.410 ;
        RECT 2484.190 1597.320 2507.270 1598.410 ;
        RECT 2508.110 1597.320 2531.190 1598.410 ;
        RECT 2532.030 1597.320 2555.110 1598.410 ;
        RECT 2555.950 1597.320 2579.030 1598.410 ;
        RECT 2579.870 1597.320 2599.830 1598.410 ;
        RECT 0.090 2.680 2599.830 1597.320 ;
        RECT 0.090 1.630 31.550 2.680 ;
        RECT 32.390 1.630 55.930 2.680 ;
        RECT 56.770 1.630 80.310 2.680 ;
        RECT 81.150 1.630 104.690 2.680 ;
        RECT 105.530 1.630 129.070 2.680 ;
        RECT 129.910 1.630 153.450 2.680 ;
        RECT 154.290 1.630 177.830 2.680 ;
        RECT 178.670 1.630 202.210 2.680 ;
        RECT 203.050 1.630 226.590 2.680 ;
        RECT 227.430 1.630 250.970 2.680 ;
        RECT 251.810 1.630 275.350 2.680 ;
        RECT 276.190 1.630 299.730 2.680 ;
        RECT 300.570 1.630 324.110 2.680 ;
        RECT 324.950 1.630 348.490 2.680 ;
        RECT 349.330 1.630 372.870 2.680 ;
        RECT 373.710 1.630 397.250 2.680 ;
        RECT 398.090 1.630 421.630 2.680 ;
        RECT 422.470 1.630 446.010 2.680 ;
        RECT 446.850 1.630 470.390 2.680 ;
        RECT 471.230 1.630 494.770 2.680 ;
        RECT 495.610 1.630 519.150 2.680 ;
        RECT 519.990 1.630 543.530 2.680 ;
        RECT 544.370 1.630 567.910 2.680 ;
        RECT 568.750 1.630 592.290 2.680 ;
        RECT 593.130 1.630 616.670 2.680 ;
        RECT 617.510 1.630 641.050 2.680 ;
        RECT 641.890 1.630 665.430 2.680 ;
        RECT 666.270 1.630 689.810 2.680 ;
        RECT 690.650 1.630 714.190 2.680 ;
        RECT 715.030 1.630 738.570 2.680 ;
        RECT 739.410 1.630 762.950 2.680 ;
        RECT 763.790 1.630 787.330 2.680 ;
        RECT 788.170 1.630 811.710 2.680 ;
        RECT 812.550 1.630 836.090 2.680 ;
        RECT 836.930 1.630 860.470 2.680 ;
        RECT 861.310 1.630 884.850 2.680 ;
        RECT 885.690 1.630 909.230 2.680 ;
        RECT 910.070 1.630 933.610 2.680 ;
        RECT 934.450 1.630 957.990 2.680 ;
        RECT 958.830 1.630 982.370 2.680 ;
        RECT 983.210 1.630 1006.750 2.680 ;
        RECT 1007.590 1.630 1031.130 2.680 ;
        RECT 1031.970 1.630 1055.510 2.680 ;
        RECT 1056.350 1.630 1079.890 2.680 ;
        RECT 1080.730 1.630 1104.270 2.680 ;
        RECT 1105.110 1.630 1128.650 2.680 ;
        RECT 1129.490 1.630 1153.030 2.680 ;
        RECT 1153.870 1.630 1177.410 2.680 ;
        RECT 1178.250 1.630 1201.790 2.680 ;
        RECT 1202.630 1.630 1226.170 2.680 ;
        RECT 1227.010 1.630 1250.550 2.680 ;
        RECT 1251.390 1.630 1274.930 2.680 ;
        RECT 1275.770 1.630 1299.310 2.680 ;
        RECT 1300.150 1.630 1323.690 2.680 ;
        RECT 1324.530 1.630 1348.070 2.680 ;
        RECT 1348.910 1.630 1372.450 2.680 ;
        RECT 1373.290 1.630 1396.830 2.680 ;
        RECT 1397.670 1.630 1421.210 2.680 ;
        RECT 1422.050 1.630 1445.590 2.680 ;
        RECT 1446.430 1.630 1469.970 2.680 ;
        RECT 1470.810 1.630 1494.350 2.680 ;
        RECT 1495.190 1.630 1518.730 2.680 ;
        RECT 1519.570 1.630 1543.110 2.680 ;
        RECT 1543.950 1.630 1567.490 2.680 ;
        RECT 1568.330 1.630 1591.870 2.680 ;
        RECT 1592.710 1.630 1616.250 2.680 ;
        RECT 1617.090 1.630 1640.630 2.680 ;
        RECT 1641.470 1.630 1665.010 2.680 ;
        RECT 1665.850 1.630 1689.390 2.680 ;
        RECT 1690.230 1.630 1713.770 2.680 ;
        RECT 1714.610 1.630 1738.150 2.680 ;
        RECT 1738.990 1.630 1762.530 2.680 ;
        RECT 1763.370 1.630 1786.910 2.680 ;
        RECT 1787.750 1.630 1811.290 2.680 ;
        RECT 1812.130 1.630 1835.670 2.680 ;
        RECT 1836.510 1.630 1860.050 2.680 ;
        RECT 1860.890 1.630 1884.430 2.680 ;
        RECT 1885.270 1.630 1908.810 2.680 ;
        RECT 1909.650 1.630 1933.190 2.680 ;
        RECT 1934.030 1.630 1957.570 2.680 ;
        RECT 1958.410 1.630 1981.950 2.680 ;
        RECT 1982.790 1.630 2006.330 2.680 ;
        RECT 2007.170 1.630 2030.710 2.680 ;
        RECT 2031.550 1.630 2055.090 2.680 ;
        RECT 2055.930 1.630 2079.470 2.680 ;
        RECT 2080.310 1.630 2103.850 2.680 ;
        RECT 2104.690 1.630 2128.230 2.680 ;
        RECT 2129.070 1.630 2152.610 2.680 ;
        RECT 2153.450 1.630 2176.990 2.680 ;
        RECT 2177.830 1.630 2201.370 2.680 ;
        RECT 2202.210 1.630 2225.750 2.680 ;
        RECT 2226.590 1.630 2250.130 2.680 ;
        RECT 2250.970 1.630 2274.510 2.680 ;
        RECT 2275.350 1.630 2298.890 2.680 ;
        RECT 2299.730 1.630 2323.270 2.680 ;
        RECT 2324.110 1.630 2347.650 2.680 ;
        RECT 2348.490 1.630 2372.030 2.680 ;
        RECT 2372.870 1.630 2396.410 2.680 ;
        RECT 2397.250 1.630 2420.790 2.680 ;
        RECT 2421.630 1.630 2445.170 2.680 ;
        RECT 2446.010 1.630 2469.550 2.680 ;
        RECT 2470.390 1.630 2493.930 2.680 ;
        RECT 2494.770 1.630 2518.310 2.680 ;
        RECT 2519.150 1.630 2542.690 2.680 ;
        RECT 2543.530 1.630 2567.070 2.680 ;
        RECT 2567.910 1.630 2599.830 2.680 ;
      LAYER met3 ;
        RECT 0.065 1531.040 2598.935 1588.645 ;
        RECT 0.065 1529.640 2597.200 1531.040 ;
        RECT 0.065 1522.880 2598.935 1529.640 ;
        RECT 0.065 1521.480 2597.200 1522.880 ;
        RECT 0.065 1514.720 2598.935 1521.480 ;
        RECT 0.065 1513.320 2597.200 1514.720 ;
        RECT 0.065 1506.560 2598.935 1513.320 ;
        RECT 0.065 1505.160 2597.200 1506.560 ;
        RECT 0.065 1498.400 2598.935 1505.160 ;
        RECT 0.065 1497.000 2597.200 1498.400 ;
        RECT 0.065 1490.240 2598.935 1497.000 ;
        RECT 2.800 1488.840 2597.200 1490.240 ;
        RECT 0.065 1482.080 2598.935 1488.840 ;
        RECT 2.800 1480.680 2597.200 1482.080 ;
        RECT 0.065 1473.920 2598.935 1480.680 ;
        RECT 2.800 1472.520 2597.200 1473.920 ;
        RECT 0.065 1465.760 2598.935 1472.520 ;
        RECT 2.800 1464.360 2597.200 1465.760 ;
        RECT 0.065 1457.600 2598.935 1464.360 ;
        RECT 2.800 1456.200 2597.200 1457.600 ;
        RECT 0.065 1449.440 2598.935 1456.200 ;
        RECT 2.800 1448.040 2597.200 1449.440 ;
        RECT 0.065 1441.280 2598.935 1448.040 ;
        RECT 2.800 1439.880 2597.200 1441.280 ;
        RECT 0.065 1433.120 2598.935 1439.880 ;
        RECT 2.800 1431.720 2597.200 1433.120 ;
        RECT 0.065 1424.960 2598.935 1431.720 ;
        RECT 2.800 1423.560 2597.200 1424.960 ;
        RECT 0.065 1416.800 2598.935 1423.560 ;
        RECT 2.800 1415.400 2597.200 1416.800 ;
        RECT 0.065 1408.640 2598.935 1415.400 ;
        RECT 2.800 1407.240 2597.200 1408.640 ;
        RECT 0.065 1400.480 2598.935 1407.240 ;
        RECT 2.800 1399.080 2597.200 1400.480 ;
        RECT 0.065 1392.320 2598.935 1399.080 ;
        RECT 2.800 1390.920 2597.200 1392.320 ;
        RECT 0.065 1384.160 2598.935 1390.920 ;
        RECT 2.800 1382.760 2597.200 1384.160 ;
        RECT 0.065 1376.000 2598.935 1382.760 ;
        RECT 2.800 1374.600 2597.200 1376.000 ;
        RECT 0.065 1367.840 2598.935 1374.600 ;
        RECT 2.800 1366.440 2597.200 1367.840 ;
        RECT 0.065 1359.680 2598.935 1366.440 ;
        RECT 2.800 1358.280 2597.200 1359.680 ;
        RECT 0.065 1351.520 2598.935 1358.280 ;
        RECT 2.800 1350.120 2597.200 1351.520 ;
        RECT 0.065 1343.360 2598.935 1350.120 ;
        RECT 2.800 1341.960 2597.200 1343.360 ;
        RECT 0.065 1335.200 2598.935 1341.960 ;
        RECT 2.800 1333.800 2597.200 1335.200 ;
        RECT 0.065 1327.040 2598.935 1333.800 ;
        RECT 2.800 1325.640 2597.200 1327.040 ;
        RECT 0.065 1318.880 2598.935 1325.640 ;
        RECT 2.800 1317.480 2597.200 1318.880 ;
        RECT 0.065 1310.720 2598.935 1317.480 ;
        RECT 2.800 1309.320 2597.200 1310.720 ;
        RECT 0.065 1302.560 2598.935 1309.320 ;
        RECT 2.800 1301.160 2597.200 1302.560 ;
        RECT 0.065 1294.400 2598.935 1301.160 ;
        RECT 2.800 1293.000 2597.200 1294.400 ;
        RECT 0.065 1286.240 2598.935 1293.000 ;
        RECT 2.800 1284.840 2597.200 1286.240 ;
        RECT 0.065 1278.080 2598.935 1284.840 ;
        RECT 2.800 1276.680 2597.200 1278.080 ;
        RECT 0.065 1269.920 2598.935 1276.680 ;
        RECT 2.800 1268.520 2597.200 1269.920 ;
        RECT 0.065 1261.760 2598.935 1268.520 ;
        RECT 2.800 1260.360 2597.200 1261.760 ;
        RECT 0.065 1253.600 2598.935 1260.360 ;
        RECT 2.800 1252.200 2597.200 1253.600 ;
        RECT 0.065 1245.440 2598.935 1252.200 ;
        RECT 2.800 1244.040 2597.200 1245.440 ;
        RECT 0.065 1237.280 2598.935 1244.040 ;
        RECT 2.800 1235.880 2597.200 1237.280 ;
        RECT 0.065 1229.120 2598.935 1235.880 ;
        RECT 2.800 1227.720 2597.200 1229.120 ;
        RECT 0.065 1220.960 2598.935 1227.720 ;
        RECT 2.800 1219.560 2597.200 1220.960 ;
        RECT 0.065 1212.800 2598.935 1219.560 ;
        RECT 2.800 1211.400 2597.200 1212.800 ;
        RECT 0.065 1204.640 2598.935 1211.400 ;
        RECT 2.800 1203.240 2597.200 1204.640 ;
        RECT 0.065 1196.480 2598.935 1203.240 ;
        RECT 2.800 1195.080 2597.200 1196.480 ;
        RECT 0.065 1188.320 2598.935 1195.080 ;
        RECT 2.800 1186.920 2597.200 1188.320 ;
        RECT 0.065 1180.160 2598.935 1186.920 ;
        RECT 2.800 1178.760 2597.200 1180.160 ;
        RECT 0.065 1172.000 2598.935 1178.760 ;
        RECT 2.800 1170.600 2597.200 1172.000 ;
        RECT 0.065 1163.840 2598.935 1170.600 ;
        RECT 2.800 1162.440 2597.200 1163.840 ;
        RECT 0.065 1155.680 2598.935 1162.440 ;
        RECT 2.800 1154.280 2597.200 1155.680 ;
        RECT 0.065 1147.520 2598.935 1154.280 ;
        RECT 2.800 1146.120 2597.200 1147.520 ;
        RECT 0.065 1139.360 2598.935 1146.120 ;
        RECT 2.800 1137.960 2597.200 1139.360 ;
        RECT 0.065 1131.200 2598.935 1137.960 ;
        RECT 2.800 1129.800 2597.200 1131.200 ;
        RECT 0.065 1123.040 2598.935 1129.800 ;
        RECT 2.800 1121.640 2597.200 1123.040 ;
        RECT 0.065 1114.880 2598.935 1121.640 ;
        RECT 2.800 1113.480 2597.200 1114.880 ;
        RECT 0.065 1106.720 2598.935 1113.480 ;
        RECT 2.800 1105.320 2597.200 1106.720 ;
        RECT 0.065 1098.560 2598.935 1105.320 ;
        RECT 2.800 1097.160 2597.200 1098.560 ;
        RECT 0.065 1090.400 2598.935 1097.160 ;
        RECT 2.800 1089.000 2597.200 1090.400 ;
        RECT 0.065 1082.240 2598.935 1089.000 ;
        RECT 2.800 1080.840 2597.200 1082.240 ;
        RECT 0.065 1074.080 2598.935 1080.840 ;
        RECT 2.800 1072.680 2597.200 1074.080 ;
        RECT 0.065 1065.920 2598.935 1072.680 ;
        RECT 2.800 1064.520 2597.200 1065.920 ;
        RECT 0.065 1057.760 2598.935 1064.520 ;
        RECT 2.800 1056.360 2597.200 1057.760 ;
        RECT 0.065 1049.600 2598.935 1056.360 ;
        RECT 2.800 1048.200 2597.200 1049.600 ;
        RECT 0.065 1041.440 2598.935 1048.200 ;
        RECT 2.800 1040.040 2597.200 1041.440 ;
        RECT 0.065 1033.280 2598.935 1040.040 ;
        RECT 2.800 1031.880 2597.200 1033.280 ;
        RECT 0.065 1025.120 2598.935 1031.880 ;
        RECT 2.800 1023.720 2597.200 1025.120 ;
        RECT 0.065 1016.960 2598.935 1023.720 ;
        RECT 2.800 1015.560 2597.200 1016.960 ;
        RECT 0.065 1008.800 2598.935 1015.560 ;
        RECT 2.800 1007.400 2597.200 1008.800 ;
        RECT 0.065 1000.640 2598.935 1007.400 ;
        RECT 2.800 999.240 2597.200 1000.640 ;
        RECT 0.065 992.480 2598.935 999.240 ;
        RECT 2.800 991.080 2597.200 992.480 ;
        RECT 0.065 984.320 2598.935 991.080 ;
        RECT 2.800 982.920 2597.200 984.320 ;
        RECT 0.065 976.160 2598.935 982.920 ;
        RECT 2.800 974.760 2597.200 976.160 ;
        RECT 0.065 968.000 2598.935 974.760 ;
        RECT 2.800 966.600 2597.200 968.000 ;
        RECT 0.065 959.840 2598.935 966.600 ;
        RECT 2.800 958.440 2597.200 959.840 ;
        RECT 0.065 951.680 2598.935 958.440 ;
        RECT 2.800 950.280 2597.200 951.680 ;
        RECT 0.065 943.520 2598.935 950.280 ;
        RECT 2.800 942.120 2597.200 943.520 ;
        RECT 0.065 935.360 2598.935 942.120 ;
        RECT 2.800 933.960 2597.200 935.360 ;
        RECT 0.065 927.200 2598.935 933.960 ;
        RECT 2.800 925.800 2597.200 927.200 ;
        RECT 0.065 919.040 2598.935 925.800 ;
        RECT 2.800 917.640 2597.200 919.040 ;
        RECT 0.065 910.880 2598.935 917.640 ;
        RECT 2.800 909.480 2597.200 910.880 ;
        RECT 0.065 902.720 2598.935 909.480 ;
        RECT 2.800 901.320 2597.200 902.720 ;
        RECT 0.065 894.560 2598.935 901.320 ;
        RECT 2.800 893.160 2597.200 894.560 ;
        RECT 0.065 886.400 2598.935 893.160 ;
        RECT 2.800 885.000 2597.200 886.400 ;
        RECT 0.065 878.240 2598.935 885.000 ;
        RECT 2.800 876.840 2597.200 878.240 ;
        RECT 0.065 870.080 2598.935 876.840 ;
        RECT 2.800 868.680 2597.200 870.080 ;
        RECT 0.065 861.920 2598.935 868.680 ;
        RECT 2.800 860.520 2597.200 861.920 ;
        RECT 0.065 853.760 2598.935 860.520 ;
        RECT 2.800 852.360 2597.200 853.760 ;
        RECT 0.065 845.600 2598.935 852.360 ;
        RECT 2.800 844.200 2597.200 845.600 ;
        RECT 0.065 837.440 2598.935 844.200 ;
        RECT 2.800 836.040 2597.200 837.440 ;
        RECT 0.065 829.280 2598.935 836.040 ;
        RECT 2.800 827.880 2597.200 829.280 ;
        RECT 0.065 821.120 2598.935 827.880 ;
        RECT 2.800 819.720 2597.200 821.120 ;
        RECT 0.065 812.960 2598.935 819.720 ;
        RECT 2.800 811.560 2597.200 812.960 ;
        RECT 0.065 804.800 2598.935 811.560 ;
        RECT 2.800 803.400 2597.200 804.800 ;
        RECT 0.065 796.640 2598.935 803.400 ;
        RECT 2.800 795.240 2597.200 796.640 ;
        RECT 0.065 788.480 2598.935 795.240 ;
        RECT 2.800 787.080 2597.200 788.480 ;
        RECT 0.065 780.320 2598.935 787.080 ;
        RECT 2.800 778.920 2597.200 780.320 ;
        RECT 0.065 772.160 2598.935 778.920 ;
        RECT 2.800 770.760 2597.200 772.160 ;
        RECT 0.065 764.000 2598.935 770.760 ;
        RECT 2.800 762.600 2597.200 764.000 ;
        RECT 0.065 755.840 2598.935 762.600 ;
        RECT 2.800 754.440 2597.200 755.840 ;
        RECT 0.065 747.680 2598.935 754.440 ;
        RECT 2.800 746.280 2597.200 747.680 ;
        RECT 0.065 739.520 2598.935 746.280 ;
        RECT 2.800 738.120 2597.200 739.520 ;
        RECT 0.065 731.360 2598.935 738.120 ;
        RECT 2.800 729.960 2597.200 731.360 ;
        RECT 0.065 723.200 2598.935 729.960 ;
        RECT 2.800 721.800 2597.200 723.200 ;
        RECT 0.065 715.040 2598.935 721.800 ;
        RECT 2.800 713.640 2597.200 715.040 ;
        RECT 0.065 706.880 2598.935 713.640 ;
        RECT 2.800 705.480 2597.200 706.880 ;
        RECT 0.065 698.720 2598.935 705.480 ;
        RECT 2.800 697.320 2597.200 698.720 ;
        RECT 0.065 690.560 2598.935 697.320 ;
        RECT 2.800 689.160 2597.200 690.560 ;
        RECT 0.065 682.400 2598.935 689.160 ;
        RECT 2.800 681.000 2597.200 682.400 ;
        RECT 0.065 674.240 2598.935 681.000 ;
        RECT 2.800 672.840 2597.200 674.240 ;
        RECT 0.065 666.080 2598.935 672.840 ;
        RECT 2.800 664.680 2597.200 666.080 ;
        RECT 0.065 657.920 2598.935 664.680 ;
        RECT 2.800 656.520 2597.200 657.920 ;
        RECT 0.065 649.760 2598.935 656.520 ;
        RECT 2.800 648.360 2597.200 649.760 ;
        RECT 0.065 641.600 2598.935 648.360 ;
        RECT 2.800 640.200 2597.200 641.600 ;
        RECT 0.065 633.440 2598.935 640.200 ;
        RECT 2.800 632.040 2597.200 633.440 ;
        RECT 0.065 625.280 2598.935 632.040 ;
        RECT 2.800 623.880 2597.200 625.280 ;
        RECT 0.065 617.120 2598.935 623.880 ;
        RECT 2.800 615.720 2597.200 617.120 ;
        RECT 0.065 608.960 2598.935 615.720 ;
        RECT 2.800 607.560 2597.200 608.960 ;
        RECT 0.065 600.800 2598.935 607.560 ;
        RECT 2.800 599.400 2597.200 600.800 ;
        RECT 0.065 592.640 2598.935 599.400 ;
        RECT 2.800 591.240 2597.200 592.640 ;
        RECT 0.065 584.480 2598.935 591.240 ;
        RECT 2.800 583.080 2597.200 584.480 ;
        RECT 0.065 576.320 2598.935 583.080 ;
        RECT 2.800 574.920 2597.200 576.320 ;
        RECT 0.065 568.160 2598.935 574.920 ;
        RECT 2.800 566.760 2597.200 568.160 ;
        RECT 0.065 560.000 2598.935 566.760 ;
        RECT 2.800 558.600 2597.200 560.000 ;
        RECT 0.065 551.840 2598.935 558.600 ;
        RECT 2.800 550.440 2597.200 551.840 ;
        RECT 0.065 543.680 2598.935 550.440 ;
        RECT 2.800 542.280 2597.200 543.680 ;
        RECT 0.065 535.520 2598.935 542.280 ;
        RECT 2.800 534.120 2597.200 535.520 ;
        RECT 0.065 527.360 2598.935 534.120 ;
        RECT 2.800 525.960 2597.200 527.360 ;
        RECT 0.065 519.200 2598.935 525.960 ;
        RECT 2.800 517.800 2597.200 519.200 ;
        RECT 0.065 511.040 2598.935 517.800 ;
        RECT 2.800 509.640 2597.200 511.040 ;
        RECT 0.065 502.880 2598.935 509.640 ;
        RECT 2.800 501.480 2597.200 502.880 ;
        RECT 0.065 494.720 2598.935 501.480 ;
        RECT 2.800 493.320 2597.200 494.720 ;
        RECT 0.065 486.560 2598.935 493.320 ;
        RECT 2.800 485.160 2597.200 486.560 ;
        RECT 0.065 478.400 2598.935 485.160 ;
        RECT 2.800 477.000 2597.200 478.400 ;
        RECT 0.065 470.240 2598.935 477.000 ;
        RECT 2.800 468.840 2597.200 470.240 ;
        RECT 0.065 462.080 2598.935 468.840 ;
        RECT 2.800 460.680 2597.200 462.080 ;
        RECT 0.065 453.920 2598.935 460.680 ;
        RECT 2.800 452.520 2597.200 453.920 ;
        RECT 0.065 445.760 2598.935 452.520 ;
        RECT 2.800 444.360 2597.200 445.760 ;
        RECT 0.065 437.600 2598.935 444.360 ;
        RECT 2.800 436.200 2597.200 437.600 ;
        RECT 0.065 429.440 2598.935 436.200 ;
        RECT 2.800 428.040 2597.200 429.440 ;
        RECT 0.065 421.280 2598.935 428.040 ;
        RECT 2.800 419.880 2597.200 421.280 ;
        RECT 0.065 413.120 2598.935 419.880 ;
        RECT 2.800 411.720 2597.200 413.120 ;
        RECT 0.065 404.960 2598.935 411.720 ;
        RECT 2.800 403.560 2597.200 404.960 ;
        RECT 0.065 396.800 2598.935 403.560 ;
        RECT 2.800 395.400 2597.200 396.800 ;
        RECT 0.065 388.640 2598.935 395.400 ;
        RECT 2.800 387.240 2597.200 388.640 ;
        RECT 0.065 380.480 2598.935 387.240 ;
        RECT 2.800 379.080 2597.200 380.480 ;
        RECT 0.065 372.320 2598.935 379.080 ;
        RECT 2.800 370.920 2597.200 372.320 ;
        RECT 0.065 364.160 2598.935 370.920 ;
        RECT 2.800 362.760 2597.200 364.160 ;
        RECT 0.065 356.000 2598.935 362.760 ;
        RECT 2.800 354.600 2597.200 356.000 ;
        RECT 0.065 347.840 2598.935 354.600 ;
        RECT 2.800 346.440 2597.200 347.840 ;
        RECT 0.065 339.680 2598.935 346.440 ;
        RECT 2.800 338.280 2597.200 339.680 ;
        RECT 0.065 331.520 2598.935 338.280 ;
        RECT 2.800 330.120 2597.200 331.520 ;
        RECT 0.065 323.360 2598.935 330.120 ;
        RECT 2.800 321.960 2597.200 323.360 ;
        RECT 0.065 315.200 2598.935 321.960 ;
        RECT 2.800 313.800 2597.200 315.200 ;
        RECT 0.065 307.040 2598.935 313.800 ;
        RECT 2.800 305.640 2597.200 307.040 ;
        RECT 0.065 298.880 2598.935 305.640 ;
        RECT 2.800 297.480 2597.200 298.880 ;
        RECT 0.065 290.720 2598.935 297.480 ;
        RECT 2.800 289.320 2597.200 290.720 ;
        RECT 0.065 282.560 2598.935 289.320 ;
        RECT 2.800 281.160 2597.200 282.560 ;
        RECT 0.065 274.400 2598.935 281.160 ;
        RECT 2.800 273.000 2597.200 274.400 ;
        RECT 0.065 266.240 2598.935 273.000 ;
        RECT 2.800 264.840 2597.200 266.240 ;
        RECT 0.065 258.080 2598.935 264.840 ;
        RECT 2.800 256.680 2597.200 258.080 ;
        RECT 0.065 249.920 2598.935 256.680 ;
        RECT 2.800 248.520 2597.200 249.920 ;
        RECT 0.065 241.760 2598.935 248.520 ;
        RECT 2.800 240.360 2597.200 241.760 ;
        RECT 0.065 233.600 2598.935 240.360 ;
        RECT 2.800 232.200 2597.200 233.600 ;
        RECT 0.065 225.440 2598.935 232.200 ;
        RECT 2.800 224.040 2597.200 225.440 ;
        RECT 0.065 217.280 2598.935 224.040 ;
        RECT 2.800 215.880 2597.200 217.280 ;
        RECT 0.065 209.120 2598.935 215.880 ;
        RECT 2.800 207.720 2597.200 209.120 ;
        RECT 0.065 200.960 2598.935 207.720 ;
        RECT 2.800 199.560 2597.200 200.960 ;
        RECT 0.065 192.800 2598.935 199.560 ;
        RECT 2.800 191.400 2597.200 192.800 ;
        RECT 0.065 184.640 2598.935 191.400 ;
        RECT 2.800 183.240 2597.200 184.640 ;
        RECT 0.065 176.480 2598.935 183.240 ;
        RECT 2.800 175.080 2597.200 176.480 ;
        RECT 0.065 168.320 2598.935 175.080 ;
        RECT 2.800 166.920 2597.200 168.320 ;
        RECT 0.065 160.160 2598.935 166.920 ;
        RECT 2.800 158.760 2597.200 160.160 ;
        RECT 0.065 152.000 2598.935 158.760 ;
        RECT 2.800 150.600 2597.200 152.000 ;
        RECT 0.065 143.840 2598.935 150.600 ;
        RECT 2.800 142.440 2597.200 143.840 ;
        RECT 0.065 135.680 2598.935 142.440 ;
        RECT 2.800 134.280 2597.200 135.680 ;
        RECT 0.065 127.520 2598.935 134.280 ;
        RECT 2.800 126.120 2597.200 127.520 ;
        RECT 0.065 119.360 2598.935 126.120 ;
        RECT 2.800 117.960 2597.200 119.360 ;
        RECT 0.065 111.200 2598.935 117.960 ;
        RECT 2.800 109.800 2597.200 111.200 ;
        RECT 0.065 103.040 2598.935 109.800 ;
        RECT 0.065 101.640 2597.200 103.040 ;
        RECT 0.065 94.880 2598.935 101.640 ;
        RECT 0.065 93.480 2597.200 94.880 ;
        RECT 0.065 86.720 2598.935 93.480 ;
        RECT 0.065 85.320 2597.200 86.720 ;
        RECT 0.065 78.560 2598.935 85.320 ;
        RECT 0.065 77.160 2597.200 78.560 ;
        RECT 0.065 70.400 2598.935 77.160 ;
        RECT 0.065 69.000 2597.200 70.400 ;
        RECT 0.065 10.715 2598.935 69.000 ;
      LAYER met4 ;
        RECT 17.775 104.895 48.570 1414.905 ;
        RECT 52.470 104.895 53.670 1414.905 ;
        RECT 57.570 1046.220 88.570 1414.905 ;
        RECT 92.470 1046.220 93.670 1414.905 ;
        RECT 97.570 1046.220 128.570 1414.905 ;
        RECT 132.470 1046.220 133.670 1414.905 ;
        RECT 137.570 1046.220 168.570 1414.905 ;
        RECT 172.470 1046.220 173.670 1414.905 ;
        RECT 177.570 1046.220 208.570 1414.905 ;
        RECT 212.470 1046.220 213.670 1414.905 ;
        RECT 217.570 1046.220 248.570 1414.905 ;
        RECT 252.470 1046.840 253.670 1414.905 ;
        RECT 257.570 1046.840 288.570 1414.905 ;
        RECT 252.470 1046.560 288.570 1046.840 ;
        RECT 292.470 1046.560 293.670 1414.905 ;
        RECT 252.470 1046.220 293.670 1046.560 ;
        RECT 297.570 1046.560 328.570 1414.905 ;
        RECT 332.470 1046.560 333.670 1414.905 ;
        RECT 297.570 1046.220 333.670 1046.560 ;
        RECT 337.570 1046.220 368.570 1414.905 ;
        RECT 372.470 1046.220 373.670 1414.905 ;
        RECT 377.570 1046.220 408.570 1414.905 ;
        RECT 412.470 1046.220 413.670 1414.905 ;
        RECT 417.570 1046.220 448.570 1414.905 ;
        RECT 452.470 1046.840 453.670 1414.905 ;
        RECT 457.570 1046.840 488.570 1414.905 ;
        RECT 452.470 1046.220 488.570 1046.840 ;
        RECT 492.470 1046.220 493.670 1414.905 ;
        RECT 497.570 1046.560 528.570 1414.905 ;
        RECT 532.470 1046.560 533.670 1414.905 ;
        RECT 497.570 1046.220 533.670 1046.560 ;
        RECT 537.570 1046.220 568.570 1414.905 ;
        RECT 572.470 1046.220 573.670 1414.905 ;
        RECT 577.570 1046.220 608.570 1414.905 ;
        RECT 612.470 1046.840 613.670 1414.905 ;
        RECT 617.570 1046.840 648.570 1414.905 ;
        RECT 612.470 1046.220 648.570 1046.840 ;
        RECT 652.470 1046.220 653.670 1414.905 ;
        RECT 657.570 1046.560 688.570 1414.905 ;
        RECT 692.470 1046.560 693.670 1414.905 ;
        RECT 657.570 1046.220 693.670 1046.560 ;
        RECT 697.570 1046.220 728.570 1414.905 ;
        RECT 732.470 1046.220 733.670 1414.905 ;
        RECT 737.570 1046.220 768.570 1414.905 ;
        RECT 772.470 1046.220 773.670 1414.905 ;
        RECT 777.570 1046.220 808.570 1414.905 ;
        RECT 57.570 610.320 808.570 1046.220 ;
        RECT 57.570 104.895 88.570 610.320 ;
        RECT 92.470 104.895 93.670 610.320 ;
        RECT 97.570 104.895 128.570 610.320 ;
        RECT 132.470 104.895 133.670 610.320 ;
        RECT 137.570 104.895 168.570 610.320 ;
        RECT 172.470 104.895 173.670 610.320 ;
        RECT 177.570 609.920 373.670 610.320 ;
        RECT 177.570 609.700 213.670 609.920 ;
        RECT 177.570 104.895 208.570 609.700 ;
        RECT 212.470 104.895 213.670 609.700 ;
        RECT 217.570 609.700 253.670 609.920 ;
        RECT 217.570 104.895 248.570 609.700 ;
        RECT 252.470 104.895 253.670 609.700 ;
        RECT 257.570 609.700 293.670 609.920 ;
        RECT 257.570 104.895 288.570 609.700 ;
        RECT 292.470 104.895 293.670 609.700 ;
        RECT 297.570 609.700 333.670 609.920 ;
        RECT 297.570 104.895 328.570 609.700 ;
        RECT 332.470 104.895 333.670 609.700 ;
        RECT 337.570 609.700 373.670 609.920 ;
        RECT 337.570 104.895 368.570 609.700 ;
        RECT 372.470 104.895 373.670 609.700 ;
        RECT 377.570 104.895 408.570 610.320 ;
        RECT 412.470 609.920 448.570 610.320 ;
        RECT 412.470 104.895 413.670 609.920 ;
        RECT 417.570 104.895 448.570 609.920 ;
        RECT 452.470 609.920 493.670 610.320 ;
        RECT 452.470 104.895 453.670 609.920 ;
        RECT 457.570 609.700 493.670 609.920 ;
        RECT 457.570 104.895 488.570 609.700 ;
        RECT 492.470 104.895 493.670 609.700 ;
        RECT 497.570 609.700 533.670 610.320 ;
        RECT 497.570 104.895 528.570 609.700 ;
        RECT 532.470 104.895 533.670 609.700 ;
        RECT 537.570 104.895 568.570 610.320 ;
        RECT 572.470 104.895 573.670 610.320 ;
        RECT 577.570 104.895 608.570 610.320 ;
        RECT 612.470 609.920 648.570 610.320 ;
        RECT 612.470 104.895 613.670 609.920 ;
        RECT 617.570 104.895 648.570 609.920 ;
        RECT 652.470 104.895 653.670 610.320 ;
        RECT 657.570 104.895 688.570 610.320 ;
        RECT 692.470 104.895 693.670 610.320 ;
        RECT 697.570 104.895 728.570 610.320 ;
        RECT 732.470 104.895 733.670 610.320 ;
        RECT 737.570 104.895 768.570 610.320 ;
        RECT 772.470 104.895 773.670 610.320 ;
        RECT 777.570 104.895 808.570 610.320 ;
        RECT 812.470 104.895 813.670 1414.905 ;
        RECT 817.570 104.895 848.570 1414.905 ;
        RECT 852.470 104.895 853.670 1414.905 ;
        RECT 857.570 104.895 888.570 1414.905 ;
        RECT 892.470 104.895 893.670 1414.905 ;
        RECT 897.570 104.895 928.570 1414.905 ;
        RECT 932.470 104.895 933.670 1414.905 ;
        RECT 937.570 104.895 968.570 1414.905 ;
        RECT 972.470 104.895 973.670 1414.905 ;
        RECT 977.570 104.895 1008.570 1414.905 ;
        RECT 1012.470 104.895 1013.670 1414.905 ;
        RECT 1017.570 104.895 1048.570 1414.905 ;
        RECT 1052.470 104.895 1053.670 1414.905 ;
        RECT 1057.570 104.895 1088.570 1414.905 ;
        RECT 1092.470 104.895 1093.670 1414.905 ;
        RECT 1097.570 104.895 1128.570 1414.905 ;
        RECT 1132.470 104.895 1133.670 1414.905 ;
        RECT 1137.570 104.895 1168.570 1414.905 ;
        RECT 1172.470 104.895 1173.670 1414.905 ;
        RECT 1177.570 778.540 1208.570 1414.905 ;
        RECT 1212.470 778.540 1213.670 1414.905 ;
        RECT 1177.570 769.965 1213.670 778.540 ;
        RECT 1217.570 778.540 1248.570 1414.905 ;
        RECT 1252.470 778.540 1253.670 1414.905 ;
        RECT 1217.570 769.965 1253.670 778.540 ;
        RECT 1177.570 741.555 1253.670 769.965 ;
        RECT 1177.570 694.900 1213.670 741.555 ;
        RECT 1177.570 104.895 1208.570 694.900 ;
        RECT 1212.470 104.895 1213.670 694.900 ;
        RECT 1217.570 694.900 1253.670 741.555 ;
        RECT 1217.570 104.895 1248.570 694.900 ;
        RECT 1252.470 104.895 1253.670 694.900 ;
        RECT 1257.570 104.895 1288.570 1414.905 ;
        RECT 1292.470 104.895 1293.670 1414.905 ;
        RECT 1297.570 104.895 1328.570 1414.905 ;
        RECT 1332.470 104.895 1333.670 1414.905 ;
        RECT 1337.570 104.895 1368.570 1414.905 ;
        RECT 1372.470 104.895 1373.670 1414.905 ;
        RECT 1377.570 1046.220 1408.570 1414.905 ;
        RECT 1412.470 1046.220 1413.670 1414.905 ;
        RECT 1417.570 1046.220 1448.570 1414.905 ;
        RECT 1452.470 1046.220 1453.670 1414.905 ;
        RECT 1457.570 1046.220 1488.570 1414.905 ;
        RECT 1492.470 1046.220 1493.670 1414.905 ;
        RECT 1497.570 1046.220 1528.570 1414.905 ;
        RECT 1532.470 1046.220 1533.670 1414.905 ;
        RECT 1537.570 1046.220 1568.570 1414.905 ;
        RECT 1572.470 1046.220 1573.670 1414.905 ;
        RECT 1577.570 1046.220 1608.570 1414.905 ;
        RECT 1612.470 1046.840 1613.670 1414.905 ;
        RECT 1617.570 1046.840 1648.570 1414.905 ;
        RECT 1612.470 1046.220 1648.570 1046.840 ;
        RECT 1652.470 1046.840 1653.670 1414.905 ;
        RECT 1657.570 1046.840 1688.570 1414.905 ;
        RECT 1652.470 1046.560 1688.570 1046.840 ;
        RECT 1692.470 1046.560 1693.670 1414.905 ;
        RECT 1652.470 1046.220 1693.670 1046.560 ;
        RECT 1697.570 1046.560 1728.570 1414.905 ;
        RECT 1732.470 1046.560 1733.670 1414.905 ;
        RECT 1697.570 1046.220 1733.670 1046.560 ;
        RECT 1737.570 1046.220 1768.570 1414.905 ;
        RECT 1772.470 1046.220 1773.670 1414.905 ;
        RECT 1777.570 1046.220 1808.570 1414.905 ;
        RECT 1812.470 1046.840 1813.670 1414.905 ;
        RECT 1817.570 1046.840 1848.570 1414.905 ;
        RECT 1812.470 1046.220 1848.570 1046.840 ;
        RECT 1852.470 1046.840 1853.670 1414.905 ;
        RECT 1857.570 1046.840 1888.570 1414.905 ;
        RECT 1852.470 1046.560 1888.570 1046.840 ;
        RECT 1892.470 1046.560 1893.670 1414.905 ;
        RECT 1852.470 1046.220 1893.670 1046.560 ;
        RECT 1897.570 1046.560 1928.570 1414.905 ;
        RECT 1932.470 1046.560 1933.670 1414.905 ;
        RECT 1897.570 1046.220 1933.670 1046.560 ;
        RECT 1937.570 1046.220 1968.570 1414.905 ;
        RECT 1972.470 1046.220 1973.670 1414.905 ;
        RECT 1977.570 1046.220 2008.570 1414.905 ;
        RECT 2012.470 1046.220 2013.670 1414.905 ;
        RECT 2017.570 1046.220 2048.570 1414.905 ;
        RECT 2052.470 1046.840 2053.670 1414.905 ;
        RECT 2057.570 1046.840 2088.570 1414.905 ;
        RECT 2052.470 1046.220 2088.570 1046.840 ;
        RECT 2092.470 1046.220 2093.670 1414.905 ;
        RECT 1377.570 610.320 2093.670 1046.220 ;
        RECT 1377.570 104.895 1408.570 610.320 ;
        RECT 1412.470 104.895 1413.670 610.320 ;
        RECT 1417.570 104.895 1448.570 610.320 ;
        RECT 1452.470 104.895 1453.670 610.320 ;
        RECT 1457.570 609.920 1533.670 610.320 ;
        RECT 1457.570 609.700 1493.670 609.920 ;
        RECT 1457.570 104.895 1488.570 609.700 ;
        RECT 1492.470 104.895 1493.670 609.700 ;
        RECT 1497.570 609.700 1533.670 609.920 ;
        RECT 1497.570 104.895 1528.570 609.700 ;
        RECT 1532.470 104.895 1533.670 609.700 ;
        RECT 1537.570 609.700 1573.670 610.320 ;
        RECT 1537.570 104.895 1568.570 609.700 ;
        RECT 1572.470 104.895 1573.670 609.700 ;
        RECT 1577.570 609.920 1733.670 610.320 ;
        RECT 1577.570 609.700 1613.670 609.920 ;
        RECT 1577.570 104.895 1608.570 609.700 ;
        RECT 1612.470 104.895 1613.670 609.700 ;
        RECT 1617.570 609.700 1653.670 609.920 ;
        RECT 1617.570 104.895 1648.570 609.700 ;
        RECT 1652.470 104.895 1653.670 609.700 ;
        RECT 1657.570 609.700 1693.670 609.920 ;
        RECT 1657.570 104.895 1688.570 609.700 ;
        RECT 1692.470 104.895 1693.670 609.700 ;
        RECT 1697.570 609.700 1733.670 609.920 ;
        RECT 1697.570 104.895 1728.570 609.700 ;
        RECT 1732.470 104.895 1733.670 609.700 ;
        RECT 1737.570 104.895 1768.570 610.320 ;
        RECT 1772.470 104.895 1773.670 610.320 ;
        RECT 1777.570 104.895 1808.570 610.320 ;
        RECT 1812.470 609.920 1848.570 610.320 ;
        RECT 1812.470 104.895 1813.670 609.920 ;
        RECT 1817.570 104.895 1848.570 609.920 ;
        RECT 1852.470 609.920 1893.670 610.320 ;
        RECT 1852.470 104.895 1853.670 609.920 ;
        RECT 1857.570 609.700 1893.670 609.920 ;
        RECT 1857.570 104.895 1888.570 609.700 ;
        RECT 1892.470 104.895 1893.670 609.700 ;
        RECT 1897.570 609.700 1933.670 610.320 ;
        RECT 1897.570 104.895 1928.570 609.700 ;
        RECT 1932.470 104.895 1933.670 609.700 ;
        RECT 1937.570 104.895 1968.570 610.320 ;
        RECT 1972.470 104.895 1973.670 610.320 ;
        RECT 1977.570 104.895 2008.570 610.320 ;
        RECT 2012.470 609.920 2048.570 610.320 ;
        RECT 2012.470 104.895 2013.670 609.920 ;
        RECT 2017.570 104.895 2048.570 609.920 ;
        RECT 2052.470 104.895 2053.670 610.320 ;
        RECT 2057.570 104.895 2088.570 610.320 ;
        RECT 2092.470 104.895 2093.670 610.320 ;
        RECT 2097.570 104.895 2128.570 1414.905 ;
        RECT 2132.470 104.895 2133.670 1414.905 ;
        RECT 2137.570 104.895 2168.570 1414.905 ;
        RECT 2172.470 104.895 2173.670 1414.905 ;
        RECT 2177.570 104.895 2208.570 1414.905 ;
        RECT 2212.470 104.895 2213.670 1414.905 ;
        RECT 2217.570 104.895 2248.570 1414.905 ;
        RECT 2252.470 104.895 2253.670 1414.905 ;
        RECT 2257.570 104.895 2288.570 1414.905 ;
        RECT 2292.470 104.895 2293.670 1414.905 ;
        RECT 2297.570 104.895 2328.570 1414.905 ;
        RECT 2332.470 104.895 2333.670 1414.905 ;
        RECT 2337.570 104.895 2368.570 1414.905 ;
        RECT 2372.470 104.895 2373.670 1414.905 ;
        RECT 2377.570 104.895 2408.570 1414.905 ;
        RECT 2412.470 104.895 2413.670 1414.905 ;
        RECT 2417.570 104.895 2448.570 1414.905 ;
        RECT 2452.470 104.895 2453.670 1414.905 ;
        RECT 2457.570 104.895 2488.570 1414.905 ;
        RECT 2492.470 104.895 2493.670 1414.905 ;
        RECT 2497.570 104.895 2528.570 1414.905 ;
        RECT 2532.470 104.895 2533.670 1414.905 ;
        RECT 2537.570 104.895 2568.570 1414.905 ;
        RECT 2572.470 104.895 2573.670 1414.905 ;
        RECT 2577.570 104.895 2586.745 1414.905 ;
      LAYER met5 ;
        RECT 260.940 744.130 1705.100 750.500 ;
        RECT 260.940 704.130 1705.100 732.730 ;
        RECT 260.940 664.130 1705.100 692.730 ;
        RECT 260.940 624.130 1705.100 652.730 ;
        RECT 260.940 584.130 1705.100 612.730 ;
        RECT 260.940 544.130 1705.100 572.730 ;
        RECT 260.940 504.130 1705.100 532.730 ;
        RECT 260.940 464.130 1705.100 492.730 ;
        RECT 260.940 424.130 1705.100 452.730 ;
        RECT 260.940 384.130 1705.100 412.730 ;
        RECT 260.940 344.130 1705.100 372.730 ;
        RECT 260.940 327.300 1705.100 332.730 ;
  END
END picosoc
END LIBRARY

