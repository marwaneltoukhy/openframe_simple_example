magic
tech sky130A
magscale 1 2
timestamp 1693307806
<< obsli1 >>
rect 1104 2159 518880 317713
<< obsm1 >>
rect 14 1912 519970 318368
<< metal2 >>
rect 3974 319520 4030 320000
rect 8758 319520 8814 320000
rect 13542 319520 13598 320000
rect 18326 319520 18382 320000
rect 23110 319520 23166 320000
rect 27894 319520 27950 320000
rect 32678 319520 32734 320000
rect 37462 319520 37518 320000
rect 42246 319520 42302 320000
rect 47030 319520 47086 320000
rect 51814 319520 51870 320000
rect 56598 319520 56654 320000
rect 61382 319520 61438 320000
rect 66166 319520 66222 320000
rect 70950 319520 71006 320000
rect 75734 319520 75790 320000
rect 80518 319520 80574 320000
rect 85302 319520 85358 320000
rect 90086 319520 90142 320000
rect 94870 319520 94926 320000
rect 99654 319520 99710 320000
rect 104438 319520 104494 320000
rect 109222 319520 109278 320000
rect 114006 319520 114062 320000
rect 118790 319520 118846 320000
rect 123574 319520 123630 320000
rect 128358 319520 128414 320000
rect 133142 319520 133198 320000
rect 137926 319520 137982 320000
rect 142710 319520 142766 320000
rect 147494 319520 147550 320000
rect 152278 319520 152334 320000
rect 157062 319520 157118 320000
rect 161846 319520 161902 320000
rect 166630 319520 166686 320000
rect 171414 319520 171470 320000
rect 176198 319520 176254 320000
rect 180982 319520 181038 320000
rect 185766 319520 185822 320000
rect 190550 319520 190606 320000
rect 195334 319520 195390 320000
rect 200118 319520 200174 320000
rect 204902 319520 204958 320000
rect 209686 319520 209742 320000
rect 214470 319520 214526 320000
rect 219254 319520 219310 320000
rect 224038 319520 224094 320000
rect 228822 319520 228878 320000
rect 233606 319520 233662 320000
rect 238390 319520 238446 320000
rect 243174 319520 243230 320000
rect 247958 319520 248014 320000
rect 252742 319520 252798 320000
rect 257526 319520 257582 320000
rect 262310 319520 262366 320000
rect 267094 319520 267150 320000
rect 271878 319520 271934 320000
rect 276662 319520 276718 320000
rect 281446 319520 281502 320000
rect 286230 319520 286286 320000
rect 291014 319520 291070 320000
rect 295798 319520 295854 320000
rect 300582 319520 300638 320000
rect 305366 319520 305422 320000
rect 310150 319520 310206 320000
rect 314934 319520 314990 320000
rect 319718 319520 319774 320000
rect 324502 319520 324558 320000
rect 329286 319520 329342 320000
rect 334070 319520 334126 320000
rect 338854 319520 338910 320000
rect 343638 319520 343694 320000
rect 348422 319520 348478 320000
rect 353206 319520 353262 320000
rect 357990 319520 358046 320000
rect 362774 319520 362830 320000
rect 367558 319520 367614 320000
rect 372342 319520 372398 320000
rect 377126 319520 377182 320000
rect 381910 319520 381966 320000
rect 386694 319520 386750 320000
rect 391478 319520 391534 320000
rect 396262 319520 396318 320000
rect 401046 319520 401102 320000
rect 405830 319520 405886 320000
rect 410614 319520 410670 320000
rect 415398 319520 415454 320000
rect 420182 319520 420238 320000
rect 424966 319520 425022 320000
rect 429750 319520 429806 320000
rect 434534 319520 434590 320000
rect 439318 319520 439374 320000
rect 444102 319520 444158 320000
rect 448886 319520 448942 320000
rect 453670 319520 453726 320000
rect 458454 319520 458510 320000
rect 463238 319520 463294 320000
rect 468022 319520 468078 320000
rect 472806 319520 472862 320000
rect 477590 319520 477646 320000
rect 482374 319520 482430 320000
rect 487158 319520 487214 320000
rect 491942 319520 491998 320000
rect 496726 319520 496782 320000
rect 501510 319520 501566 320000
rect 506294 319520 506350 320000
rect 511078 319520 511134 320000
rect 515862 319520 515918 320000
rect 6366 0 6422 480
rect 11242 0 11298 480
rect 16118 0 16174 480
rect 20994 0 21050 480
rect 25870 0 25926 480
rect 30746 0 30802 480
rect 35622 0 35678 480
rect 40498 0 40554 480
rect 45374 0 45430 480
rect 50250 0 50306 480
rect 55126 0 55182 480
rect 60002 0 60058 480
rect 64878 0 64934 480
rect 69754 0 69810 480
rect 74630 0 74686 480
rect 79506 0 79562 480
rect 84382 0 84438 480
rect 89258 0 89314 480
rect 94134 0 94190 480
rect 99010 0 99066 480
rect 103886 0 103942 480
rect 108762 0 108818 480
rect 113638 0 113694 480
rect 118514 0 118570 480
rect 123390 0 123446 480
rect 128266 0 128322 480
rect 133142 0 133198 480
rect 138018 0 138074 480
rect 142894 0 142950 480
rect 147770 0 147826 480
rect 152646 0 152702 480
rect 157522 0 157578 480
rect 162398 0 162454 480
rect 167274 0 167330 480
rect 172150 0 172206 480
rect 177026 0 177082 480
rect 181902 0 181958 480
rect 186778 0 186834 480
rect 191654 0 191710 480
rect 196530 0 196586 480
rect 201406 0 201462 480
rect 206282 0 206338 480
rect 211158 0 211214 480
rect 216034 0 216090 480
rect 220910 0 220966 480
rect 225786 0 225842 480
rect 230662 0 230718 480
rect 235538 0 235594 480
rect 240414 0 240470 480
rect 245290 0 245346 480
rect 250166 0 250222 480
rect 255042 0 255098 480
rect 259918 0 259974 480
rect 264794 0 264850 480
rect 269670 0 269726 480
rect 274546 0 274602 480
rect 279422 0 279478 480
rect 284298 0 284354 480
rect 289174 0 289230 480
rect 294050 0 294106 480
rect 298926 0 298982 480
rect 303802 0 303858 480
rect 308678 0 308734 480
rect 313554 0 313610 480
rect 318430 0 318486 480
rect 323306 0 323362 480
rect 328182 0 328238 480
rect 333058 0 333114 480
rect 337934 0 337990 480
rect 342810 0 342866 480
rect 347686 0 347742 480
rect 352562 0 352618 480
rect 357438 0 357494 480
rect 362314 0 362370 480
rect 367190 0 367246 480
rect 372066 0 372122 480
rect 376942 0 376998 480
rect 381818 0 381874 480
rect 386694 0 386750 480
rect 391570 0 391626 480
rect 396446 0 396502 480
rect 401322 0 401378 480
rect 406198 0 406254 480
rect 411074 0 411130 480
rect 415950 0 416006 480
rect 420826 0 420882 480
rect 425702 0 425758 480
rect 430578 0 430634 480
rect 435454 0 435510 480
rect 440330 0 440386 480
rect 445206 0 445262 480
rect 450082 0 450138 480
rect 454958 0 455014 480
rect 459834 0 459890 480
rect 464710 0 464766 480
rect 469586 0 469642 480
rect 474462 0 474518 480
rect 479338 0 479394 480
rect 484214 0 484270 480
rect 489090 0 489146 480
rect 493966 0 494022 480
rect 498842 0 498898 480
rect 503718 0 503774 480
rect 508594 0 508650 480
rect 513470 0 513526 480
<< obsm2 >>
rect 18 319464 3918 319682
rect 4086 319464 8702 319682
rect 8870 319464 13486 319682
rect 13654 319464 18270 319682
rect 18438 319464 23054 319682
rect 23222 319464 27838 319682
rect 28006 319464 32622 319682
rect 32790 319464 37406 319682
rect 37574 319464 42190 319682
rect 42358 319464 46974 319682
rect 47142 319464 51758 319682
rect 51926 319464 56542 319682
rect 56710 319464 61326 319682
rect 61494 319464 66110 319682
rect 66278 319464 70894 319682
rect 71062 319464 75678 319682
rect 75846 319464 80462 319682
rect 80630 319464 85246 319682
rect 85414 319464 90030 319682
rect 90198 319464 94814 319682
rect 94982 319464 99598 319682
rect 99766 319464 104382 319682
rect 104550 319464 109166 319682
rect 109334 319464 113950 319682
rect 114118 319464 118734 319682
rect 118902 319464 123518 319682
rect 123686 319464 128302 319682
rect 128470 319464 133086 319682
rect 133254 319464 137870 319682
rect 138038 319464 142654 319682
rect 142822 319464 147438 319682
rect 147606 319464 152222 319682
rect 152390 319464 157006 319682
rect 157174 319464 161790 319682
rect 161958 319464 166574 319682
rect 166742 319464 171358 319682
rect 171526 319464 176142 319682
rect 176310 319464 180926 319682
rect 181094 319464 185710 319682
rect 185878 319464 190494 319682
rect 190662 319464 195278 319682
rect 195446 319464 200062 319682
rect 200230 319464 204846 319682
rect 205014 319464 209630 319682
rect 209798 319464 214414 319682
rect 214582 319464 219198 319682
rect 219366 319464 223982 319682
rect 224150 319464 228766 319682
rect 228934 319464 233550 319682
rect 233718 319464 238334 319682
rect 238502 319464 243118 319682
rect 243286 319464 247902 319682
rect 248070 319464 252686 319682
rect 252854 319464 257470 319682
rect 257638 319464 262254 319682
rect 262422 319464 267038 319682
rect 267206 319464 271822 319682
rect 271990 319464 276606 319682
rect 276774 319464 281390 319682
rect 281558 319464 286174 319682
rect 286342 319464 290958 319682
rect 291126 319464 295742 319682
rect 295910 319464 300526 319682
rect 300694 319464 305310 319682
rect 305478 319464 310094 319682
rect 310262 319464 314878 319682
rect 315046 319464 319662 319682
rect 319830 319464 324446 319682
rect 324614 319464 329230 319682
rect 329398 319464 334014 319682
rect 334182 319464 338798 319682
rect 338966 319464 343582 319682
rect 343750 319464 348366 319682
rect 348534 319464 353150 319682
rect 353318 319464 357934 319682
rect 358102 319464 362718 319682
rect 362886 319464 367502 319682
rect 367670 319464 372286 319682
rect 372454 319464 377070 319682
rect 377238 319464 381854 319682
rect 382022 319464 386638 319682
rect 386806 319464 391422 319682
rect 391590 319464 396206 319682
rect 396374 319464 400990 319682
rect 401158 319464 405774 319682
rect 405942 319464 410558 319682
rect 410726 319464 415342 319682
rect 415510 319464 420126 319682
rect 420294 319464 424910 319682
rect 425078 319464 429694 319682
rect 429862 319464 434478 319682
rect 434646 319464 439262 319682
rect 439430 319464 444046 319682
rect 444214 319464 448830 319682
rect 448998 319464 453614 319682
rect 453782 319464 458398 319682
rect 458566 319464 463182 319682
rect 463350 319464 467966 319682
rect 468134 319464 472750 319682
rect 472918 319464 477534 319682
rect 477702 319464 482318 319682
rect 482486 319464 487102 319682
rect 487270 319464 491886 319682
rect 492054 319464 496670 319682
rect 496838 319464 501454 319682
rect 501622 319464 506238 319682
rect 506406 319464 511022 319682
rect 511190 319464 515806 319682
rect 515974 319464 519966 319682
rect 18 536 519966 319464
rect 18 326 6310 536
rect 6478 326 11186 536
rect 11354 326 16062 536
rect 16230 326 20938 536
rect 21106 326 25814 536
rect 25982 326 30690 536
rect 30858 326 35566 536
rect 35734 326 40442 536
rect 40610 326 45318 536
rect 45486 326 50194 536
rect 50362 326 55070 536
rect 55238 326 59946 536
rect 60114 326 64822 536
rect 64990 326 69698 536
rect 69866 326 74574 536
rect 74742 326 79450 536
rect 79618 326 84326 536
rect 84494 326 89202 536
rect 89370 326 94078 536
rect 94246 326 98954 536
rect 99122 326 103830 536
rect 103998 326 108706 536
rect 108874 326 113582 536
rect 113750 326 118458 536
rect 118626 326 123334 536
rect 123502 326 128210 536
rect 128378 326 133086 536
rect 133254 326 137962 536
rect 138130 326 142838 536
rect 143006 326 147714 536
rect 147882 326 152590 536
rect 152758 326 157466 536
rect 157634 326 162342 536
rect 162510 326 167218 536
rect 167386 326 172094 536
rect 172262 326 176970 536
rect 177138 326 181846 536
rect 182014 326 186722 536
rect 186890 326 191598 536
rect 191766 326 196474 536
rect 196642 326 201350 536
rect 201518 326 206226 536
rect 206394 326 211102 536
rect 211270 326 215978 536
rect 216146 326 220854 536
rect 221022 326 225730 536
rect 225898 326 230606 536
rect 230774 326 235482 536
rect 235650 326 240358 536
rect 240526 326 245234 536
rect 245402 326 250110 536
rect 250278 326 254986 536
rect 255154 326 259862 536
rect 260030 326 264738 536
rect 264906 326 269614 536
rect 269782 326 274490 536
rect 274658 326 279366 536
rect 279534 326 284242 536
rect 284410 326 289118 536
rect 289286 326 293994 536
rect 294162 326 298870 536
rect 299038 326 303746 536
rect 303914 326 308622 536
rect 308790 326 313498 536
rect 313666 326 318374 536
rect 318542 326 323250 536
rect 323418 326 328126 536
rect 328294 326 333002 536
rect 333170 326 337878 536
rect 338046 326 342754 536
rect 342922 326 347630 536
rect 347798 326 352506 536
rect 352674 326 357382 536
rect 357550 326 362258 536
rect 362426 326 367134 536
rect 367302 326 372010 536
rect 372178 326 376886 536
rect 377054 326 381762 536
rect 381930 326 386638 536
rect 386806 326 391514 536
rect 391682 326 396390 536
rect 396558 326 401266 536
rect 401434 326 406142 536
rect 406310 326 411018 536
rect 411186 326 415894 536
rect 416062 326 420770 536
rect 420938 326 425646 536
rect 425814 326 430522 536
rect 430690 326 435398 536
rect 435566 326 440274 536
rect 440442 326 445150 536
rect 445318 326 450026 536
rect 450194 326 454902 536
rect 455070 326 459778 536
rect 459946 326 464654 536
rect 464822 326 469530 536
rect 469698 326 474406 536
rect 474574 326 479282 536
rect 479450 326 484158 536
rect 484326 326 489034 536
rect 489202 326 493910 536
rect 494078 326 498786 536
rect 498954 326 503662 536
rect 503830 326 508538 536
rect 508706 326 513414 536
rect 513582 326 519966 536
<< metal3 >>
rect 519520 306008 520000 306128
rect 519520 304376 520000 304496
rect 519520 302744 520000 302864
rect 519520 301112 520000 301232
rect 519520 299480 520000 299600
rect 0 297848 480 297968
rect 519520 297848 520000 297968
rect 0 296216 480 296336
rect 519520 296216 520000 296336
rect 0 294584 480 294704
rect 519520 294584 520000 294704
rect 0 292952 480 293072
rect 519520 292952 520000 293072
rect 0 291320 480 291440
rect 519520 291320 520000 291440
rect 0 289688 480 289808
rect 519520 289688 520000 289808
rect 0 288056 480 288176
rect 519520 288056 520000 288176
rect 0 286424 480 286544
rect 519520 286424 520000 286544
rect 0 284792 480 284912
rect 519520 284792 520000 284912
rect 0 283160 480 283280
rect 519520 283160 520000 283280
rect 0 281528 480 281648
rect 519520 281528 520000 281648
rect 0 279896 480 280016
rect 519520 279896 520000 280016
rect 0 278264 480 278384
rect 519520 278264 520000 278384
rect 0 276632 480 276752
rect 519520 276632 520000 276752
rect 0 275000 480 275120
rect 519520 275000 520000 275120
rect 0 273368 480 273488
rect 519520 273368 520000 273488
rect 0 271736 480 271856
rect 519520 271736 520000 271856
rect 0 270104 480 270224
rect 519520 270104 520000 270224
rect 0 268472 480 268592
rect 519520 268472 520000 268592
rect 0 266840 480 266960
rect 519520 266840 520000 266960
rect 0 265208 480 265328
rect 519520 265208 520000 265328
rect 0 263576 480 263696
rect 519520 263576 520000 263696
rect 0 261944 480 262064
rect 519520 261944 520000 262064
rect 0 260312 480 260432
rect 519520 260312 520000 260432
rect 0 258680 480 258800
rect 519520 258680 520000 258800
rect 0 257048 480 257168
rect 519520 257048 520000 257168
rect 0 255416 480 255536
rect 519520 255416 520000 255536
rect 0 253784 480 253904
rect 519520 253784 520000 253904
rect 0 252152 480 252272
rect 519520 252152 520000 252272
rect 0 250520 480 250640
rect 519520 250520 520000 250640
rect 0 248888 480 249008
rect 519520 248888 520000 249008
rect 0 247256 480 247376
rect 519520 247256 520000 247376
rect 0 245624 480 245744
rect 519520 245624 520000 245744
rect 0 243992 480 244112
rect 519520 243992 520000 244112
rect 0 242360 480 242480
rect 519520 242360 520000 242480
rect 0 240728 480 240848
rect 519520 240728 520000 240848
rect 0 239096 480 239216
rect 519520 239096 520000 239216
rect 0 237464 480 237584
rect 519520 237464 520000 237584
rect 0 235832 480 235952
rect 519520 235832 520000 235952
rect 0 234200 480 234320
rect 519520 234200 520000 234320
rect 0 232568 480 232688
rect 519520 232568 520000 232688
rect 0 230936 480 231056
rect 519520 230936 520000 231056
rect 0 229304 480 229424
rect 519520 229304 520000 229424
rect 0 227672 480 227792
rect 519520 227672 520000 227792
rect 0 226040 480 226160
rect 519520 226040 520000 226160
rect 0 224408 480 224528
rect 519520 224408 520000 224528
rect 0 222776 480 222896
rect 519520 222776 520000 222896
rect 0 221144 480 221264
rect 519520 221144 520000 221264
rect 0 219512 480 219632
rect 519520 219512 520000 219632
rect 0 217880 480 218000
rect 519520 217880 520000 218000
rect 0 216248 480 216368
rect 519520 216248 520000 216368
rect 0 214616 480 214736
rect 519520 214616 520000 214736
rect 0 212984 480 213104
rect 519520 212984 520000 213104
rect 0 211352 480 211472
rect 519520 211352 520000 211472
rect 0 209720 480 209840
rect 519520 209720 520000 209840
rect 0 208088 480 208208
rect 519520 208088 520000 208208
rect 0 206456 480 206576
rect 519520 206456 520000 206576
rect 0 204824 480 204944
rect 519520 204824 520000 204944
rect 0 203192 480 203312
rect 519520 203192 520000 203312
rect 0 201560 480 201680
rect 519520 201560 520000 201680
rect 0 199928 480 200048
rect 519520 199928 520000 200048
rect 0 198296 480 198416
rect 519520 198296 520000 198416
rect 0 196664 480 196784
rect 519520 196664 520000 196784
rect 0 195032 480 195152
rect 519520 195032 520000 195152
rect 0 193400 480 193520
rect 519520 193400 520000 193520
rect 0 191768 480 191888
rect 519520 191768 520000 191888
rect 0 190136 480 190256
rect 519520 190136 520000 190256
rect 0 188504 480 188624
rect 519520 188504 520000 188624
rect 0 186872 480 186992
rect 519520 186872 520000 186992
rect 0 185240 480 185360
rect 519520 185240 520000 185360
rect 0 183608 480 183728
rect 519520 183608 520000 183728
rect 0 181976 480 182096
rect 519520 181976 520000 182096
rect 0 180344 480 180464
rect 519520 180344 520000 180464
rect 0 178712 480 178832
rect 519520 178712 520000 178832
rect 0 177080 480 177200
rect 519520 177080 520000 177200
rect 0 175448 480 175568
rect 519520 175448 520000 175568
rect 0 173816 480 173936
rect 519520 173816 520000 173936
rect 0 172184 480 172304
rect 519520 172184 520000 172304
rect 0 170552 480 170672
rect 519520 170552 520000 170672
rect 0 168920 480 169040
rect 519520 168920 520000 169040
rect 0 167288 480 167408
rect 519520 167288 520000 167408
rect 0 165656 480 165776
rect 519520 165656 520000 165776
rect 0 164024 480 164144
rect 519520 164024 520000 164144
rect 0 162392 480 162512
rect 519520 162392 520000 162512
rect 0 160760 480 160880
rect 519520 160760 520000 160880
rect 0 159128 480 159248
rect 519520 159128 520000 159248
rect 0 157496 480 157616
rect 519520 157496 520000 157616
rect 0 155864 480 155984
rect 519520 155864 520000 155984
rect 0 154232 480 154352
rect 519520 154232 520000 154352
rect 0 152600 480 152720
rect 519520 152600 520000 152720
rect 0 150968 480 151088
rect 519520 150968 520000 151088
rect 0 149336 480 149456
rect 519520 149336 520000 149456
rect 0 147704 480 147824
rect 519520 147704 520000 147824
rect 0 146072 480 146192
rect 519520 146072 520000 146192
rect 0 144440 480 144560
rect 519520 144440 520000 144560
rect 0 142808 480 142928
rect 519520 142808 520000 142928
rect 0 141176 480 141296
rect 519520 141176 520000 141296
rect 0 139544 480 139664
rect 519520 139544 520000 139664
rect 0 137912 480 138032
rect 519520 137912 520000 138032
rect 0 136280 480 136400
rect 519520 136280 520000 136400
rect 0 134648 480 134768
rect 519520 134648 520000 134768
rect 0 133016 480 133136
rect 519520 133016 520000 133136
rect 0 131384 480 131504
rect 519520 131384 520000 131504
rect 0 129752 480 129872
rect 519520 129752 520000 129872
rect 0 128120 480 128240
rect 519520 128120 520000 128240
rect 0 126488 480 126608
rect 519520 126488 520000 126608
rect 0 124856 480 124976
rect 519520 124856 520000 124976
rect 0 123224 480 123344
rect 519520 123224 520000 123344
rect 0 121592 480 121712
rect 519520 121592 520000 121712
rect 0 119960 480 120080
rect 519520 119960 520000 120080
rect 0 118328 480 118448
rect 519520 118328 520000 118448
rect 0 116696 480 116816
rect 519520 116696 520000 116816
rect 0 115064 480 115184
rect 519520 115064 520000 115184
rect 0 113432 480 113552
rect 519520 113432 520000 113552
rect 0 111800 480 111920
rect 519520 111800 520000 111920
rect 0 110168 480 110288
rect 519520 110168 520000 110288
rect 0 108536 480 108656
rect 519520 108536 520000 108656
rect 0 106904 480 107024
rect 519520 106904 520000 107024
rect 0 105272 480 105392
rect 519520 105272 520000 105392
rect 0 103640 480 103760
rect 519520 103640 520000 103760
rect 0 102008 480 102128
rect 519520 102008 520000 102128
rect 0 100376 480 100496
rect 519520 100376 520000 100496
rect 0 98744 480 98864
rect 519520 98744 520000 98864
rect 0 97112 480 97232
rect 519520 97112 520000 97232
rect 0 95480 480 95600
rect 519520 95480 520000 95600
rect 0 93848 480 93968
rect 519520 93848 520000 93968
rect 0 92216 480 92336
rect 519520 92216 520000 92336
rect 0 90584 480 90704
rect 519520 90584 520000 90704
rect 0 88952 480 89072
rect 519520 88952 520000 89072
rect 0 87320 480 87440
rect 519520 87320 520000 87440
rect 0 85688 480 85808
rect 519520 85688 520000 85808
rect 0 84056 480 84176
rect 519520 84056 520000 84176
rect 0 82424 480 82544
rect 519520 82424 520000 82544
rect 0 80792 480 80912
rect 519520 80792 520000 80912
rect 0 79160 480 79280
rect 519520 79160 520000 79280
rect 0 77528 480 77648
rect 519520 77528 520000 77648
rect 0 75896 480 76016
rect 519520 75896 520000 76016
rect 0 74264 480 74384
rect 519520 74264 520000 74384
rect 0 72632 480 72752
rect 519520 72632 520000 72752
rect 0 71000 480 71120
rect 519520 71000 520000 71120
rect 0 69368 480 69488
rect 519520 69368 520000 69488
rect 0 67736 480 67856
rect 519520 67736 520000 67856
rect 0 66104 480 66224
rect 519520 66104 520000 66224
rect 0 64472 480 64592
rect 519520 64472 520000 64592
rect 0 62840 480 62960
rect 519520 62840 520000 62960
rect 0 61208 480 61328
rect 519520 61208 520000 61328
rect 0 59576 480 59696
rect 519520 59576 520000 59696
rect 0 57944 480 58064
rect 519520 57944 520000 58064
rect 0 56312 480 56432
rect 519520 56312 520000 56432
rect 0 54680 480 54800
rect 519520 54680 520000 54800
rect 0 53048 480 53168
rect 519520 53048 520000 53168
rect 0 51416 480 51536
rect 519520 51416 520000 51536
rect 0 49784 480 49904
rect 519520 49784 520000 49904
rect 0 48152 480 48272
rect 519520 48152 520000 48272
rect 0 46520 480 46640
rect 519520 46520 520000 46640
rect 0 44888 480 45008
rect 519520 44888 520000 45008
rect 0 43256 480 43376
rect 519520 43256 520000 43376
rect 0 41624 480 41744
rect 519520 41624 520000 41744
rect 0 39992 480 40112
rect 519520 39992 520000 40112
rect 0 38360 480 38480
rect 519520 38360 520000 38480
rect 0 36728 480 36848
rect 519520 36728 520000 36848
rect 0 35096 480 35216
rect 519520 35096 520000 35216
rect 0 33464 480 33584
rect 519520 33464 520000 33584
rect 0 31832 480 31952
rect 519520 31832 520000 31952
rect 0 30200 480 30320
rect 519520 30200 520000 30320
rect 0 28568 480 28688
rect 519520 28568 520000 28688
rect 0 26936 480 27056
rect 519520 26936 520000 27056
rect 0 25304 480 25424
rect 519520 25304 520000 25424
rect 0 23672 480 23792
rect 519520 23672 520000 23792
rect 0 22040 480 22160
rect 519520 22040 520000 22160
rect 519520 20408 520000 20528
rect 519520 18776 520000 18896
rect 519520 17144 520000 17264
rect 519520 15512 520000 15632
rect 519520 13880 520000 14000
<< obsm3 >>
rect 13 306208 519787 317729
rect 13 305928 519440 306208
rect 13 304576 519787 305928
rect 13 304296 519440 304576
rect 13 302944 519787 304296
rect 13 302664 519440 302944
rect 13 301312 519787 302664
rect 13 301032 519440 301312
rect 13 299680 519787 301032
rect 13 299400 519440 299680
rect 13 298048 519787 299400
rect 560 297768 519440 298048
rect 13 296416 519787 297768
rect 560 296136 519440 296416
rect 13 294784 519787 296136
rect 560 294504 519440 294784
rect 13 293152 519787 294504
rect 560 292872 519440 293152
rect 13 291520 519787 292872
rect 560 291240 519440 291520
rect 13 289888 519787 291240
rect 560 289608 519440 289888
rect 13 288256 519787 289608
rect 560 287976 519440 288256
rect 13 286624 519787 287976
rect 560 286344 519440 286624
rect 13 284992 519787 286344
rect 560 284712 519440 284992
rect 13 283360 519787 284712
rect 560 283080 519440 283360
rect 13 281728 519787 283080
rect 560 281448 519440 281728
rect 13 280096 519787 281448
rect 560 279816 519440 280096
rect 13 278464 519787 279816
rect 560 278184 519440 278464
rect 13 276832 519787 278184
rect 560 276552 519440 276832
rect 13 275200 519787 276552
rect 560 274920 519440 275200
rect 13 273568 519787 274920
rect 560 273288 519440 273568
rect 13 271936 519787 273288
rect 560 271656 519440 271936
rect 13 270304 519787 271656
rect 560 270024 519440 270304
rect 13 268672 519787 270024
rect 560 268392 519440 268672
rect 13 267040 519787 268392
rect 560 266760 519440 267040
rect 13 265408 519787 266760
rect 560 265128 519440 265408
rect 13 263776 519787 265128
rect 560 263496 519440 263776
rect 13 262144 519787 263496
rect 560 261864 519440 262144
rect 13 260512 519787 261864
rect 560 260232 519440 260512
rect 13 258880 519787 260232
rect 560 258600 519440 258880
rect 13 257248 519787 258600
rect 560 256968 519440 257248
rect 13 255616 519787 256968
rect 560 255336 519440 255616
rect 13 253984 519787 255336
rect 560 253704 519440 253984
rect 13 252352 519787 253704
rect 560 252072 519440 252352
rect 13 250720 519787 252072
rect 560 250440 519440 250720
rect 13 249088 519787 250440
rect 560 248808 519440 249088
rect 13 247456 519787 248808
rect 560 247176 519440 247456
rect 13 245824 519787 247176
rect 560 245544 519440 245824
rect 13 244192 519787 245544
rect 560 243912 519440 244192
rect 13 242560 519787 243912
rect 560 242280 519440 242560
rect 13 240928 519787 242280
rect 560 240648 519440 240928
rect 13 239296 519787 240648
rect 560 239016 519440 239296
rect 13 237664 519787 239016
rect 560 237384 519440 237664
rect 13 236032 519787 237384
rect 560 235752 519440 236032
rect 13 234400 519787 235752
rect 560 234120 519440 234400
rect 13 232768 519787 234120
rect 560 232488 519440 232768
rect 13 231136 519787 232488
rect 560 230856 519440 231136
rect 13 229504 519787 230856
rect 560 229224 519440 229504
rect 13 227872 519787 229224
rect 560 227592 519440 227872
rect 13 226240 519787 227592
rect 560 225960 519440 226240
rect 13 224608 519787 225960
rect 560 224328 519440 224608
rect 13 222976 519787 224328
rect 560 222696 519440 222976
rect 13 221344 519787 222696
rect 560 221064 519440 221344
rect 13 219712 519787 221064
rect 560 219432 519440 219712
rect 13 218080 519787 219432
rect 560 217800 519440 218080
rect 13 216448 519787 217800
rect 560 216168 519440 216448
rect 13 214816 519787 216168
rect 560 214536 519440 214816
rect 13 213184 519787 214536
rect 560 212904 519440 213184
rect 13 211552 519787 212904
rect 560 211272 519440 211552
rect 13 209920 519787 211272
rect 560 209640 519440 209920
rect 13 208288 519787 209640
rect 560 208008 519440 208288
rect 13 206656 519787 208008
rect 560 206376 519440 206656
rect 13 205024 519787 206376
rect 560 204744 519440 205024
rect 13 203392 519787 204744
rect 560 203112 519440 203392
rect 13 201760 519787 203112
rect 560 201480 519440 201760
rect 13 200128 519787 201480
rect 560 199848 519440 200128
rect 13 198496 519787 199848
rect 560 198216 519440 198496
rect 13 196864 519787 198216
rect 560 196584 519440 196864
rect 13 195232 519787 196584
rect 560 194952 519440 195232
rect 13 193600 519787 194952
rect 560 193320 519440 193600
rect 13 191968 519787 193320
rect 560 191688 519440 191968
rect 13 190336 519787 191688
rect 560 190056 519440 190336
rect 13 188704 519787 190056
rect 560 188424 519440 188704
rect 13 187072 519787 188424
rect 560 186792 519440 187072
rect 13 185440 519787 186792
rect 560 185160 519440 185440
rect 13 183808 519787 185160
rect 560 183528 519440 183808
rect 13 182176 519787 183528
rect 560 181896 519440 182176
rect 13 180544 519787 181896
rect 560 180264 519440 180544
rect 13 178912 519787 180264
rect 560 178632 519440 178912
rect 13 177280 519787 178632
rect 560 177000 519440 177280
rect 13 175648 519787 177000
rect 560 175368 519440 175648
rect 13 174016 519787 175368
rect 560 173736 519440 174016
rect 13 172384 519787 173736
rect 560 172104 519440 172384
rect 13 170752 519787 172104
rect 560 170472 519440 170752
rect 13 169120 519787 170472
rect 560 168840 519440 169120
rect 13 167488 519787 168840
rect 560 167208 519440 167488
rect 13 165856 519787 167208
rect 560 165576 519440 165856
rect 13 164224 519787 165576
rect 560 163944 519440 164224
rect 13 162592 519787 163944
rect 560 162312 519440 162592
rect 13 160960 519787 162312
rect 560 160680 519440 160960
rect 13 159328 519787 160680
rect 560 159048 519440 159328
rect 13 157696 519787 159048
rect 560 157416 519440 157696
rect 13 156064 519787 157416
rect 560 155784 519440 156064
rect 13 154432 519787 155784
rect 560 154152 519440 154432
rect 13 152800 519787 154152
rect 560 152520 519440 152800
rect 13 151168 519787 152520
rect 560 150888 519440 151168
rect 13 149536 519787 150888
rect 560 149256 519440 149536
rect 13 147904 519787 149256
rect 560 147624 519440 147904
rect 13 146272 519787 147624
rect 560 145992 519440 146272
rect 13 144640 519787 145992
rect 560 144360 519440 144640
rect 13 143008 519787 144360
rect 560 142728 519440 143008
rect 13 141376 519787 142728
rect 560 141096 519440 141376
rect 13 139744 519787 141096
rect 560 139464 519440 139744
rect 13 138112 519787 139464
rect 560 137832 519440 138112
rect 13 136480 519787 137832
rect 560 136200 519440 136480
rect 13 134848 519787 136200
rect 560 134568 519440 134848
rect 13 133216 519787 134568
rect 560 132936 519440 133216
rect 13 131584 519787 132936
rect 560 131304 519440 131584
rect 13 129952 519787 131304
rect 560 129672 519440 129952
rect 13 128320 519787 129672
rect 560 128040 519440 128320
rect 13 126688 519787 128040
rect 560 126408 519440 126688
rect 13 125056 519787 126408
rect 560 124776 519440 125056
rect 13 123424 519787 124776
rect 560 123144 519440 123424
rect 13 121792 519787 123144
rect 560 121512 519440 121792
rect 13 120160 519787 121512
rect 560 119880 519440 120160
rect 13 118528 519787 119880
rect 560 118248 519440 118528
rect 13 116896 519787 118248
rect 560 116616 519440 116896
rect 13 115264 519787 116616
rect 560 114984 519440 115264
rect 13 113632 519787 114984
rect 560 113352 519440 113632
rect 13 112000 519787 113352
rect 560 111720 519440 112000
rect 13 110368 519787 111720
rect 560 110088 519440 110368
rect 13 108736 519787 110088
rect 560 108456 519440 108736
rect 13 107104 519787 108456
rect 560 106824 519440 107104
rect 13 105472 519787 106824
rect 560 105192 519440 105472
rect 13 103840 519787 105192
rect 560 103560 519440 103840
rect 13 102208 519787 103560
rect 560 101928 519440 102208
rect 13 100576 519787 101928
rect 560 100296 519440 100576
rect 13 98944 519787 100296
rect 560 98664 519440 98944
rect 13 97312 519787 98664
rect 560 97032 519440 97312
rect 13 95680 519787 97032
rect 560 95400 519440 95680
rect 13 94048 519787 95400
rect 560 93768 519440 94048
rect 13 92416 519787 93768
rect 560 92136 519440 92416
rect 13 90784 519787 92136
rect 560 90504 519440 90784
rect 13 89152 519787 90504
rect 560 88872 519440 89152
rect 13 87520 519787 88872
rect 560 87240 519440 87520
rect 13 85888 519787 87240
rect 560 85608 519440 85888
rect 13 84256 519787 85608
rect 560 83976 519440 84256
rect 13 82624 519787 83976
rect 560 82344 519440 82624
rect 13 80992 519787 82344
rect 560 80712 519440 80992
rect 13 79360 519787 80712
rect 560 79080 519440 79360
rect 13 77728 519787 79080
rect 560 77448 519440 77728
rect 13 76096 519787 77448
rect 560 75816 519440 76096
rect 13 74464 519787 75816
rect 560 74184 519440 74464
rect 13 72832 519787 74184
rect 560 72552 519440 72832
rect 13 71200 519787 72552
rect 560 70920 519440 71200
rect 13 69568 519787 70920
rect 560 69288 519440 69568
rect 13 67936 519787 69288
rect 560 67656 519440 67936
rect 13 66304 519787 67656
rect 560 66024 519440 66304
rect 13 64672 519787 66024
rect 560 64392 519440 64672
rect 13 63040 519787 64392
rect 560 62760 519440 63040
rect 13 61408 519787 62760
rect 560 61128 519440 61408
rect 13 59776 519787 61128
rect 560 59496 519440 59776
rect 13 58144 519787 59496
rect 560 57864 519440 58144
rect 13 56512 519787 57864
rect 560 56232 519440 56512
rect 13 54880 519787 56232
rect 560 54600 519440 54880
rect 13 53248 519787 54600
rect 560 52968 519440 53248
rect 13 51616 519787 52968
rect 560 51336 519440 51616
rect 13 49984 519787 51336
rect 560 49704 519440 49984
rect 13 48352 519787 49704
rect 560 48072 519440 48352
rect 13 46720 519787 48072
rect 560 46440 519440 46720
rect 13 45088 519787 46440
rect 560 44808 519440 45088
rect 13 43456 519787 44808
rect 560 43176 519440 43456
rect 13 41824 519787 43176
rect 560 41544 519440 41824
rect 13 40192 519787 41544
rect 560 39912 519440 40192
rect 13 38560 519787 39912
rect 560 38280 519440 38560
rect 13 36928 519787 38280
rect 560 36648 519440 36928
rect 13 35296 519787 36648
rect 560 35016 519440 35296
rect 13 33664 519787 35016
rect 560 33384 519440 33664
rect 13 32032 519787 33384
rect 560 31752 519440 32032
rect 13 30400 519787 31752
rect 560 30120 519440 30400
rect 13 28768 519787 30120
rect 560 28488 519440 28768
rect 13 27136 519787 28488
rect 560 26856 519440 27136
rect 13 25504 519787 26856
rect 560 25224 519440 25504
rect 13 23872 519787 25224
rect 560 23592 519440 23872
rect 13 22240 519787 23592
rect 560 21960 519440 22240
rect 13 20608 519787 21960
rect 13 20328 519440 20608
rect 13 18976 519787 20328
rect 13 18696 519440 18976
rect 13 17344 519787 18696
rect 13 17064 519440 17344
rect 13 15712 519787 17064
rect 13 15432 519440 15712
rect 13 14080 519787 15432
rect 13 13800 519440 14080
rect 13 2143 519787 13800
<< metal4 >>
rect 1794 2128 2414 317744
rect 2814 2128 3434 317744
rect 9794 2128 10414 317744
rect 10814 2128 11434 317744
rect 17794 209324 18414 317744
rect 18814 209324 19434 317744
rect 25794 209324 26414 317744
rect 26814 209324 27434 317744
rect 33794 209324 34414 317744
rect 34814 209324 35434 317744
rect 41794 209324 42414 317744
rect 42814 209324 43434 317744
rect 49794 209324 50414 317744
rect 50814 209448 51434 317744
rect 57794 209392 58414 317744
rect 58814 209324 59434 317744
rect 65794 209392 66414 317744
rect 66814 209324 67434 317744
rect 73794 209324 74414 317744
rect 74814 209324 75434 317744
rect 81794 209324 82414 317744
rect 82814 209324 83434 317744
rect 89794 209324 90414 317744
rect 90814 209448 91434 317744
rect 97794 209324 98414 317744
rect 98814 209324 99434 317744
rect 105794 209392 106414 317744
rect 106814 209324 107434 317744
rect 113794 209324 114414 317744
rect 114814 209324 115434 317744
rect 121794 209324 122414 317744
rect 122814 209448 123434 317744
rect 129794 209324 130414 317744
rect 130814 209324 131434 317744
rect 137794 209392 138414 317744
rect 138814 209324 139434 317744
rect 145794 209324 146414 317744
rect 146814 209324 147434 317744
rect 153794 209324 154414 317744
rect 154814 209324 155434 317744
rect 17794 2128 18414 121984
rect 18814 2128 19434 121984
rect 25794 2128 26414 121984
rect 26814 2128 27434 121984
rect 33794 2128 34414 121984
rect 34814 2128 35434 121984
rect 41794 2128 42414 121860
rect 42814 2128 43434 121904
rect 49794 2128 50414 121860
rect 50814 2128 51434 121904
rect 57794 2128 58414 121860
rect 58814 2128 59434 121904
rect 65794 2128 66414 121860
rect 66814 2128 67434 121904
rect 73794 2128 74414 121860
rect 74814 2128 75434 121984
rect 81794 2128 82414 121984
rect 82814 2128 83434 121904
rect 89794 2128 90414 121984
rect 90814 2128 91434 121904
rect 97794 2128 98414 121860
rect 98814 2128 99434 121984
rect 105794 2128 106414 121860
rect 106814 2128 107434 121984
rect 113794 2128 114414 121984
rect 114814 2128 115434 121984
rect 121794 2128 122414 121984
rect 122814 2128 123434 121904
rect 129794 2128 130414 121984
rect 130814 2128 131434 121984
rect 137794 2128 138414 121984
rect 138814 2128 139434 121984
rect 145794 2128 146414 121984
rect 146814 2128 147434 121984
rect 153794 2128 154414 121984
rect 154814 2128 155434 121984
rect 161794 2128 162414 317744
rect 162814 2128 163434 317744
rect 169794 2128 170414 317744
rect 170814 2128 171434 317744
rect 177794 2128 178414 317744
rect 178814 2128 179434 317744
rect 185794 2128 186414 317744
rect 186814 2128 187434 317744
rect 193794 2128 194414 317744
rect 194814 2128 195434 317744
rect 201794 2128 202414 317744
rect 202814 2128 203434 317744
rect 209794 2128 210414 317744
rect 210814 2128 211434 317744
rect 217794 2128 218414 317744
rect 218814 2128 219434 317744
rect 225794 2128 226414 317744
rect 226814 2128 227434 317744
rect 233794 2128 234414 317744
rect 234814 2128 235434 317744
rect 241794 155788 242414 317744
rect 242814 154073 243434 317744
rect 249794 155788 250414 317744
rect 241794 2128 242414 138900
rect 242814 2128 243434 148231
rect 249794 2128 250414 138900
rect 250814 2128 251434 317744
rect 257794 2128 258414 317744
rect 258814 2128 259434 317744
rect 265794 2128 266414 317744
rect 266814 2128 267434 317744
rect 273794 2128 274414 317744
rect 274814 2128 275434 317744
rect 281794 209324 282414 317744
rect 282814 209324 283434 317744
rect 289794 209324 290414 317744
rect 290814 209324 291434 317744
rect 297794 209324 298414 317744
rect 298814 209324 299434 317744
rect 305794 209324 306414 317744
rect 306814 209324 307434 317744
rect 313794 209324 314414 317744
rect 314814 209324 315434 317744
rect 321794 209324 322414 317744
rect 322814 209448 323434 317744
rect 329794 209324 330414 317744
rect 330814 209448 331434 317744
rect 337794 209392 338414 317744
rect 338814 209324 339434 317744
rect 345794 209392 346414 317744
rect 346814 209324 347434 317744
rect 353794 209324 354414 317744
rect 354814 209324 355434 317744
rect 361794 209324 362414 317744
rect 362814 209448 363434 317744
rect 369794 209324 370414 317744
rect 370814 209448 371434 317744
rect 377794 209392 378414 317744
rect 378814 209324 379434 317744
rect 385794 209392 386414 317744
rect 386814 209324 387434 317744
rect 393794 209324 394414 317744
rect 394814 209324 395434 317744
rect 401794 209324 402414 317744
rect 402814 209324 403434 317744
rect 409794 209324 410414 317744
rect 410814 209448 411434 317744
rect 417794 209324 418414 317744
rect 281794 2128 282414 121984
rect 282814 2128 283434 121984
rect 289794 2128 290414 121984
rect 290814 2128 291434 121984
rect 297794 2128 298414 121860
rect 298814 2128 299434 121904
rect 305794 2128 306414 121860
rect 306814 2128 307434 121984
rect 313794 2128 314414 121860
rect 314814 2128 315434 121984
rect 321794 2128 322414 121860
rect 322814 2128 323434 121904
rect 329794 2128 330414 121860
rect 330814 2128 331434 121904
rect 337794 2128 338414 121860
rect 338814 2128 339434 121904
rect 345794 2128 346414 121860
rect 346814 2128 347434 121984
rect 353794 2128 354414 121984
rect 354814 2128 355434 121984
rect 361794 2128 362414 121984
rect 362814 2128 363434 121904
rect 369794 2128 370414 121984
rect 370814 2128 371434 121904
rect 377794 2128 378414 121860
rect 378814 2128 379434 121984
rect 385794 2128 386414 121860
rect 386814 2128 387434 121984
rect 393794 2128 394414 121984
rect 394814 2128 395434 121984
rect 401794 2128 402414 121984
rect 402814 2128 403434 121904
rect 409794 2128 410414 121984
rect 410814 2128 411434 121984
rect 417794 2128 418414 121984
rect 418814 2128 419434 317744
rect 425794 2128 426414 317744
rect 426814 2128 427434 317744
rect 433794 2128 434414 317744
rect 434814 2128 435434 317744
rect 441794 2128 442414 317744
rect 442814 2128 443434 317744
rect 449794 2128 450414 317744
rect 450814 2128 451434 317744
rect 457794 2128 458414 317744
rect 458814 2128 459434 317744
rect 465794 2128 466414 317744
rect 466814 2128 467434 317744
rect 473794 2128 474414 317744
rect 474814 2128 475434 317744
rect 481794 2128 482414 317744
rect 482814 2128 483434 317744
rect 489794 2128 490414 317744
rect 490814 2128 491434 317744
rect 497794 2128 498414 317744
rect 498814 2128 499434 317744
rect 505794 2128 506414 317744
rect 506814 2128 507434 317744
rect 513794 2128 514414 317744
rect 514814 2128 515434 317744
<< obsm4 >>
rect 3555 20979 9714 282981
rect 10494 20979 10734 282981
rect 11514 209244 17714 282981
rect 18494 209244 18734 282981
rect 19514 209244 25714 282981
rect 26494 209244 26734 282981
rect 27514 209244 33714 282981
rect 34494 209244 34734 282981
rect 35514 209244 41714 282981
rect 42494 209244 42734 282981
rect 43514 209244 49714 282981
rect 50494 209368 50734 282981
rect 51514 209368 57714 282981
rect 50494 209312 57714 209368
rect 58494 209312 58734 282981
rect 50494 209244 58734 209312
rect 59514 209312 65714 282981
rect 66494 209312 66734 282981
rect 59514 209244 66734 209312
rect 67514 209244 73714 282981
rect 74494 209244 74734 282981
rect 75514 209244 81714 282981
rect 82494 209244 82734 282981
rect 83514 209244 89714 282981
rect 90494 209368 90734 282981
rect 91514 209368 97714 282981
rect 90494 209244 97714 209368
rect 98494 209244 98734 282981
rect 99514 209312 105714 282981
rect 106494 209312 106734 282981
rect 99514 209244 106734 209312
rect 107514 209244 113714 282981
rect 114494 209244 114734 282981
rect 115514 209244 121714 282981
rect 122494 209368 122734 282981
rect 123514 209368 129714 282981
rect 122494 209244 129714 209368
rect 130494 209244 130734 282981
rect 131514 209312 137714 282981
rect 138494 209312 138734 282981
rect 131514 209244 138734 209312
rect 139514 209244 145714 282981
rect 146494 209244 146734 282981
rect 147514 209244 153714 282981
rect 154494 209244 154734 282981
rect 155514 209244 161714 282981
rect 11514 122064 161714 209244
rect 11514 20979 17714 122064
rect 18494 20979 18734 122064
rect 19514 20979 25714 122064
rect 26494 20979 26734 122064
rect 27514 20979 33714 122064
rect 34494 20979 34734 122064
rect 35514 121984 74734 122064
rect 35514 121940 42734 121984
rect 35514 20979 41714 121940
rect 42494 20979 42734 121940
rect 43514 121940 50734 121984
rect 43514 20979 49714 121940
rect 50494 20979 50734 121940
rect 51514 121940 58734 121984
rect 51514 20979 57714 121940
rect 58494 20979 58734 121940
rect 59514 121940 66734 121984
rect 59514 20979 65714 121940
rect 66494 20979 66734 121940
rect 67514 121940 74734 121984
rect 67514 20979 73714 121940
rect 74494 20979 74734 121940
rect 75514 20979 81714 122064
rect 82494 121984 89714 122064
rect 90494 121984 98734 122064
rect 82494 20979 82734 121984
rect 83514 20979 89714 121984
rect 90494 20979 90734 121984
rect 91514 121940 98734 121984
rect 91514 20979 97714 121940
rect 98494 20979 98734 121940
rect 99514 121940 106734 122064
rect 99514 20979 105714 121940
rect 106494 20979 106734 121940
rect 107514 20979 113714 122064
rect 114494 20979 114734 122064
rect 115514 20979 121714 122064
rect 122494 121984 129714 122064
rect 122494 20979 122734 121984
rect 123514 20979 129714 121984
rect 130494 20979 130734 122064
rect 131514 20979 137714 122064
rect 138494 20979 138734 122064
rect 139514 20979 145714 122064
rect 146494 20979 146734 122064
rect 147514 20979 153714 122064
rect 154494 20979 154734 122064
rect 155514 20979 161714 122064
rect 162494 20979 162734 282981
rect 163514 20979 169714 282981
rect 170494 20979 170734 282981
rect 171514 20979 177714 282981
rect 178494 20979 178734 282981
rect 179514 20979 185714 282981
rect 186494 20979 186734 282981
rect 187514 20979 193714 282981
rect 194494 20979 194734 282981
rect 195514 20979 201714 282981
rect 202494 20979 202734 282981
rect 203514 20979 209714 282981
rect 210494 20979 210734 282981
rect 211514 20979 217714 282981
rect 218494 20979 218734 282981
rect 219514 20979 225714 282981
rect 226494 20979 226734 282981
rect 227514 20979 233714 282981
rect 234494 20979 234734 282981
rect 235514 155708 241714 282981
rect 242494 155708 242734 282981
rect 235514 153993 242734 155708
rect 243514 155708 249714 282981
rect 250494 155708 250734 282981
rect 243514 153993 250734 155708
rect 235514 148311 250734 153993
rect 235514 138980 242734 148311
rect 235514 20979 241714 138980
rect 242494 20979 242734 138980
rect 243514 138980 250734 148311
rect 243514 20979 249714 138980
rect 250494 20979 250734 138980
rect 251514 20979 257714 282981
rect 258494 20979 258734 282981
rect 259514 20979 265714 282981
rect 266494 20979 266734 282981
rect 267514 20979 273714 282981
rect 274494 20979 274734 282981
rect 275514 209244 281714 282981
rect 282494 209244 282734 282981
rect 283514 209244 289714 282981
rect 290494 209244 290734 282981
rect 291514 209244 297714 282981
rect 298494 209244 298734 282981
rect 299514 209244 305714 282981
rect 306494 209244 306734 282981
rect 307514 209244 313714 282981
rect 314494 209244 314734 282981
rect 315514 209244 321714 282981
rect 322494 209368 322734 282981
rect 323514 209368 329714 282981
rect 322494 209244 329714 209368
rect 330494 209368 330734 282981
rect 331514 209368 337714 282981
rect 330494 209312 337714 209368
rect 338494 209312 338734 282981
rect 330494 209244 338734 209312
rect 339514 209312 345714 282981
rect 346494 209312 346734 282981
rect 339514 209244 346734 209312
rect 347514 209244 353714 282981
rect 354494 209244 354734 282981
rect 355514 209244 361714 282981
rect 362494 209368 362734 282981
rect 363514 209368 369714 282981
rect 362494 209244 369714 209368
rect 370494 209368 370734 282981
rect 371514 209368 377714 282981
rect 370494 209312 377714 209368
rect 378494 209312 378734 282981
rect 370494 209244 378734 209312
rect 379514 209312 385714 282981
rect 386494 209312 386734 282981
rect 379514 209244 386734 209312
rect 387514 209244 393714 282981
rect 394494 209244 394734 282981
rect 395514 209244 401714 282981
rect 402494 209244 402734 282981
rect 403514 209244 409714 282981
rect 410494 209368 410734 282981
rect 411514 209368 417714 282981
rect 410494 209244 417714 209368
rect 418494 209244 418734 282981
rect 275514 122064 418734 209244
rect 275514 20979 281714 122064
rect 282494 20979 282734 122064
rect 283514 20979 289714 122064
rect 290494 20979 290734 122064
rect 291514 121984 306734 122064
rect 291514 121940 298734 121984
rect 291514 20979 297714 121940
rect 298494 20979 298734 121940
rect 299514 121940 306734 121984
rect 299514 20979 305714 121940
rect 306494 20979 306734 121940
rect 307514 121940 314734 122064
rect 315514 121984 346734 122064
rect 307514 20979 313714 121940
rect 314494 20979 314734 121940
rect 315514 121940 322734 121984
rect 315514 20979 321714 121940
rect 322494 20979 322734 121940
rect 323514 121940 330734 121984
rect 323514 20979 329714 121940
rect 330494 20979 330734 121940
rect 331514 121940 338734 121984
rect 331514 20979 337714 121940
rect 338494 20979 338734 121940
rect 339514 121940 346734 121984
rect 339514 20979 345714 121940
rect 346494 20979 346734 121940
rect 347514 20979 353714 122064
rect 354494 20979 354734 122064
rect 355514 20979 361714 122064
rect 362494 121984 369714 122064
rect 370494 121984 378734 122064
rect 362494 20979 362734 121984
rect 363514 20979 369714 121984
rect 370494 20979 370734 121984
rect 371514 121940 378734 121984
rect 371514 20979 377714 121940
rect 378494 20979 378734 121940
rect 379514 121940 386734 122064
rect 379514 20979 385714 121940
rect 386494 20979 386734 121940
rect 387514 20979 393714 122064
rect 394494 20979 394734 122064
rect 395514 20979 401714 122064
rect 402494 121984 409714 122064
rect 402494 20979 402734 121984
rect 403514 20979 409714 121984
rect 410494 20979 410734 122064
rect 411514 20979 417714 122064
rect 418494 20979 418734 122064
rect 419514 20979 425714 282981
rect 426494 20979 426734 282981
rect 427514 20979 433714 282981
rect 434494 20979 434734 282981
rect 435514 20979 441714 282981
rect 442494 20979 442734 282981
rect 443514 20979 449714 282981
rect 450494 20979 450734 282981
rect 451514 20979 457714 282981
rect 458494 20979 458734 282981
rect 459514 20979 465714 282981
rect 466494 20979 466734 282981
rect 467514 20979 473714 282981
rect 474494 20979 474734 282981
rect 475514 20979 481714 282981
rect 482494 20979 482734 282981
rect 483514 20979 489714 282981
rect 490494 20979 490734 282981
rect 491514 20979 497714 282981
rect 498494 20979 498734 282981
rect 499514 20979 505714 282981
rect 506494 20979 506734 282981
rect 507514 20979 513714 282981
rect 514494 20979 514734 282981
rect 515514 20979 517349 282981
<< metal5 >>
rect 1056 315886 518928 316506
rect 1056 314866 518928 315486
rect 1056 307886 518928 308506
rect 1056 306866 518928 307486
rect 1056 299886 518928 300506
rect 1056 298866 518928 299486
rect 1056 291886 518928 292506
rect 1056 290866 518928 291486
rect 1056 283886 518928 284506
rect 1056 282866 518928 283486
rect 1056 275886 518928 276506
rect 1056 274866 518928 275486
rect 1056 267886 518928 268506
rect 1056 266866 518928 267486
rect 1056 259886 518928 260506
rect 1056 258866 518928 259486
rect 1056 251886 518928 252506
rect 1056 250866 518928 251486
rect 1056 243886 518928 244506
rect 1056 242866 518928 243486
rect 1056 235886 518928 236506
rect 1056 234866 518928 235486
rect 1056 227886 518928 228506
rect 1056 226866 518928 227486
rect 1056 219886 518928 220506
rect 1056 218866 518928 219486
rect 1056 211886 518928 212506
rect 1056 210866 518928 211486
rect 1056 203886 518928 204506
rect 1056 202866 518928 203486
rect 1056 195886 518928 196506
rect 1056 194866 518928 195486
rect 1056 187886 518928 188506
rect 1056 186866 518928 187486
rect 1056 179886 518928 180506
rect 1056 178866 518928 179486
rect 1056 171886 518928 172506
rect 1056 170866 518928 171486
rect 1056 163886 518928 164506
rect 1056 162866 518928 163486
rect 1056 155886 518928 156506
rect 1056 154866 518928 155486
rect 1056 147886 518928 148506
rect 1056 146866 518928 147486
rect 1056 139886 518928 140506
rect 1056 138866 518928 139486
rect 1056 131886 518928 132506
rect 1056 130866 518928 131486
rect 1056 123886 518928 124506
rect 1056 122866 518928 123486
rect 1056 115886 518928 116506
rect 1056 114866 518928 115486
rect 1056 107886 518928 108506
rect 1056 106866 518928 107486
rect 1056 99886 518928 100506
rect 1056 98866 518928 99486
rect 1056 91886 518928 92506
rect 1056 90866 518928 91486
rect 1056 83886 518928 84506
rect 1056 82866 518928 83486
rect 1056 75886 518928 76506
rect 1056 74866 518928 75486
rect 1056 67886 518928 68506
rect 1056 66866 518928 67486
rect 1056 59886 518928 60506
rect 1056 58866 518928 59486
rect 1056 51886 518928 52506
rect 1056 50866 518928 51486
rect 1056 43886 518928 44506
rect 1056 42866 518928 43486
rect 1056 35886 518928 36506
rect 1056 34866 518928 35486
rect 1056 27886 518928 28506
rect 1056 26866 518928 27486
rect 1056 19886 518928 20506
rect 1056 18866 518928 19486
rect 1056 11886 518928 12506
rect 1056 10866 518928 11486
rect 1056 3886 518928 4506
rect 1056 2866 518928 3486
<< obsm5 >>
rect 52188 148826 341020 150100
rect 52188 140826 341020 146546
rect 52188 132826 341020 138546
rect 52188 124826 341020 130546
rect 52188 116826 341020 122546
rect 52188 108826 341020 114546
rect 52188 100826 341020 106546
rect 52188 92826 341020 98546
rect 52188 84826 341020 90546
rect 52188 76826 341020 82546
rect 52188 68826 341020 74546
rect 52188 65460 341020 66546
<< labels >>
rlabel metal4 s 2814 2128 3434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10814 2128 11434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 18814 2128 19434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 18814 209324 19434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 26814 2128 27434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 26814 209324 27434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 34814 2128 35434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 34814 209324 35434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42814 2128 43434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42814 209324 43434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50814 2128 51434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50814 209448 51434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58814 2128 59434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58814 209324 59434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66814 2128 67434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 66814 209324 67434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 74814 2128 75434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 74814 209324 75434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 82814 2128 83434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 82814 209324 83434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 90814 2128 91434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 90814 209448 91434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 98814 2128 99434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 98814 209324 99434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 106814 2128 107434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 106814 209324 107434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 114814 2128 115434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 114814 209324 115434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 122814 2128 123434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 122814 209448 123434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 130814 2128 131434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 130814 209324 131434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138814 2128 139434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138814 209324 139434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146814 2128 147434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146814 209324 147434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 154814 2128 155434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 154814 209324 155434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 162814 2128 163434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 170814 2128 171434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 178814 2128 179434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 186814 2128 187434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 194814 2128 195434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 202814 2128 203434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 210814 2128 211434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218814 2128 219434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 226814 2128 227434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 234814 2128 235434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 242814 2128 243434 148231 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 242814 154073 243434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 250814 2128 251434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 258814 2128 259434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 266814 2128 267434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 274814 2128 275434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 282814 2128 283434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 282814 209324 283434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 290814 2128 291434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 290814 209324 291434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298814 2128 299434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298814 209324 299434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 306814 2128 307434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 306814 209324 307434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 314814 2128 315434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 314814 209324 315434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 322814 2128 323434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 322814 209448 323434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 330814 2128 331434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 330814 209448 331434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 338814 2128 339434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 338814 209324 339434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 346814 2128 347434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 346814 209324 347434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 354814 2128 355434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 354814 209324 355434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 362814 2128 363434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 362814 209448 363434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 370814 2128 371434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 370814 209448 371434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378814 2128 379434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378814 209324 379434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 386814 2128 387434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 386814 209324 387434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 394814 2128 395434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 394814 209324 395434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 402814 2128 403434 121904 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 402814 209324 403434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 410814 2128 411434 121984 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 410814 209448 411434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 418814 2128 419434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 426814 2128 427434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 434814 2128 435434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 442814 2128 443434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 450814 2128 451434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 458814 2128 459434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 466814 2128 467434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 474814 2128 475434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 482814 2128 483434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 490814 2128 491434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 498814 2128 499434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 506814 2128 507434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 514814 2128 515434 317744 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3886 518928 4506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11886 518928 12506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 19886 518928 20506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 27886 518928 28506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 35886 518928 36506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 43886 518928 44506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 51886 518928 52506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 59886 518928 60506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 67886 518928 68506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 75886 518928 76506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 83886 518928 84506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 91886 518928 92506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 99886 518928 100506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 107886 518928 108506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 115886 518928 116506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 123886 518928 124506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 131886 518928 132506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 139886 518928 140506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 147886 518928 148506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 155886 518928 156506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 163886 518928 164506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 171886 518928 172506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 179886 518928 180506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 187886 518928 188506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 195886 518928 196506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 203886 518928 204506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 211886 518928 212506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 219886 518928 220506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 227886 518928 228506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 235886 518928 236506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 243886 518928 244506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 251886 518928 252506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 259886 518928 260506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 267886 518928 268506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 275886 518928 276506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 283886 518928 284506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 291886 518928 292506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 299886 518928 300506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 307886 518928 308506 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 315886 518928 316506 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9794 2128 10414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 17794 2128 18414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 17794 209324 18414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25794 2128 26414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25794 209324 26414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 33794 2128 34414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 33794 209324 34414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41794 2128 42414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41794 209324 42414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 49794 2128 50414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 49794 209324 50414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 57794 2128 58414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 57794 209392 58414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65794 2128 66414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65794 209392 66414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 209324 74414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 81794 2128 82414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 81794 209324 82414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 89794 2128 90414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 89794 209324 90414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 97794 2128 98414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 97794 209324 98414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 105794 2128 106414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 105794 209392 106414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 113794 2128 114414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 113794 209324 114414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 121794 2128 122414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 121794 209324 122414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 129794 2128 130414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 129794 209324 130414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137794 2128 138414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137794 209392 138414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145794 2128 146414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 145794 209324 146414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 153794 2128 154414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 153794 209324 154414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 161794 2128 162414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 169794 2128 170414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 177794 2128 178414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 185794 2128 186414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 193794 2128 194414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 201794 2128 202414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 209794 2128 210414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217794 2128 218414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 225794 2128 226414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 233794 2128 234414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 241794 2128 242414 138900 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 241794 155788 242414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 249794 2128 250414 138900 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 249794 155788 250414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 257794 2128 258414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 265794 2128 266414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 273794 2128 274414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 281794 2128 282414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 281794 209324 282414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 289794 2128 290414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 289794 209324 290414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297794 2128 298414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297794 209324 298414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 305794 2128 306414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 305794 209324 306414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 313794 2128 314414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 313794 209324 314414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 321794 2128 322414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 321794 209324 322414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 329794 2128 330414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 329794 209324 330414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 337794 2128 338414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 337794 209392 338414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 345794 2128 346414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 345794 209392 346414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 353794 2128 354414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 353794 209324 354414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 361794 2128 362414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 361794 209324 362414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 369794 2128 370414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 369794 209324 370414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377794 2128 378414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377794 209392 378414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385794 2128 386414 121860 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385794 209392 386414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 393794 2128 394414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 393794 209324 394414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 401794 2128 402414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 401794 209324 402414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 409794 2128 410414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 409794 209324 410414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 417794 2128 418414 121984 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 417794 209324 418414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 425794 2128 426414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 433794 2128 434414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 441794 2128 442414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 449794 2128 450414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457794 2128 458414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 465794 2128 466414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 473794 2128 474414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 481794 2128 482414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 489794 2128 490414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 497794 2128 498414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 505794 2128 506414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 513794 2128 514414 317744 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2866 518928 3486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 10866 518928 11486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18866 518928 19486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 26866 518928 27486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 34866 518928 35486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 42866 518928 43486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 50866 518928 51486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 58866 518928 59486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66866 518928 67486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 74866 518928 75486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 82866 518928 83486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 90866 518928 91486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 98866 518928 99486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 106866 518928 107486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 114866 518928 115486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 122866 518928 123486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 130866 518928 131486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 138866 518928 139486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 146866 518928 147486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 154866 518928 155486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 162866 518928 163486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 170866 518928 171486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 178866 518928 179486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 186866 518928 187486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 194866 518928 195486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 202866 518928 203486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 210866 518928 211486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 218866 518928 219486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 226866 518928 227486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 234866 518928 235486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 242866 518928 243486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 250866 518928 251486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 258866 518928 259486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 266866 518928 267486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 274866 518928 275486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 282866 518928 283486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 290866 518928 291486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 298866 518928 299486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 306866 518928 307486 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 314866 518928 315486 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 519520 18776 520000 18896 6 gpio_dm0[0]
port 3 nsew signal output
rlabel metal3 s 519520 214616 520000 214736 6 gpio_dm0[10]
port 4 nsew signal output
rlabel metal3 s 519520 234200 520000 234320 6 gpio_dm0[11]
port 5 nsew signal output
rlabel metal3 s 519520 253784 520000 253904 6 gpio_dm0[12]
port 6 nsew signal output
rlabel metal3 s 519520 273368 520000 273488 6 gpio_dm0[13]
port 7 nsew signal output
rlabel metal3 s 519520 292952 520000 293072 6 gpio_dm0[14]
port 8 nsew signal output
rlabel metal2 s 501510 319520 501566 320000 6 gpio_dm0[15]
port 9 nsew signal output
rlabel metal2 s 444102 319520 444158 320000 6 gpio_dm0[16]
port 10 nsew signal output
rlabel metal2 s 386694 319520 386750 320000 6 gpio_dm0[17]
port 11 nsew signal output
rlabel metal2 s 329286 319520 329342 320000 6 gpio_dm0[18]
port 12 nsew signal output
rlabel metal2 s 271878 319520 271934 320000 6 gpio_dm0[19]
port 13 nsew signal output
rlabel metal3 s 519520 38360 520000 38480 6 gpio_dm0[1]
port 14 nsew signal output
rlabel metal2 s 214470 319520 214526 320000 6 gpio_dm0[20]
port 15 nsew signal output
rlabel metal2 s 157062 319520 157118 320000 6 gpio_dm0[21]
port 16 nsew signal output
rlabel metal2 s 99654 319520 99710 320000 6 gpio_dm0[22]
port 17 nsew signal output
rlabel metal2 s 42246 319520 42302 320000 6 gpio_dm0[23]
port 18 nsew signal output
rlabel metal3 s 0 292952 480 293072 6 gpio_dm0[24]
port 19 nsew signal output
rlabel metal3 s 0 273368 480 273488 6 gpio_dm0[25]
port 20 nsew signal output
rlabel metal3 s 0 253784 480 253904 6 gpio_dm0[26]
port 21 nsew signal output
rlabel metal3 s 0 234200 480 234320 6 gpio_dm0[27]
port 22 nsew signal output
rlabel metal3 s 0 214616 480 214736 6 gpio_dm0[28]
port 23 nsew signal output
rlabel metal3 s 0 195032 480 195152 6 gpio_dm0[29]
port 24 nsew signal output
rlabel metal3 s 519520 57944 520000 58064 6 gpio_dm0[2]
port 25 nsew signal output
rlabel metal3 s 0 175448 480 175568 6 gpio_dm0[30]
port 26 nsew signal output
rlabel metal3 s 0 155864 480 155984 6 gpio_dm0[31]
port 27 nsew signal output
rlabel metal3 s 0 136280 480 136400 6 gpio_dm0[32]
port 28 nsew signal output
rlabel metal3 s 0 116696 480 116816 6 gpio_dm0[33]
port 29 nsew signal output
rlabel metal3 s 0 97112 480 97232 6 gpio_dm0[34]
port 30 nsew signal output
rlabel metal3 s 0 77528 480 77648 6 gpio_dm0[35]
port 31 nsew signal output
rlabel metal3 s 0 57944 480 58064 6 gpio_dm0[36]
port 32 nsew signal output
rlabel metal3 s 0 38360 480 38480 6 gpio_dm0[37]
port 33 nsew signal output
rlabel metal2 s 25870 0 25926 480 6 gpio_dm0[38]
port 34 nsew signal output
rlabel metal2 s 84382 0 84438 480 6 gpio_dm0[39]
port 35 nsew signal output
rlabel metal3 s 519520 77528 520000 77648 6 gpio_dm0[3]
port 36 nsew signal output
rlabel metal2 s 142894 0 142950 480 6 gpio_dm0[40]
port 37 nsew signal output
rlabel metal2 s 201406 0 201462 480 6 gpio_dm0[41]
port 38 nsew signal output
rlabel metal2 s 259918 0 259974 480 6 gpio_dm0[42]
port 39 nsew signal output
rlabel metal2 s 318430 0 318486 480 6 gpio_dm0[43]
port 40 nsew signal output
rlabel metal3 s 519520 97112 520000 97232 6 gpio_dm0[4]
port 41 nsew signal output
rlabel metal3 s 519520 116696 520000 116816 6 gpio_dm0[5]
port 42 nsew signal output
rlabel metal3 s 519520 136280 520000 136400 6 gpio_dm0[6]
port 43 nsew signal output
rlabel metal3 s 519520 155864 520000 155984 6 gpio_dm0[7]
port 44 nsew signal output
rlabel metal3 s 519520 175448 520000 175568 6 gpio_dm0[8]
port 45 nsew signal output
rlabel metal3 s 519520 195032 520000 195152 6 gpio_dm0[9]
port 46 nsew signal output
rlabel metal3 s 519520 17144 520000 17264 6 gpio_dm1[0]
port 47 nsew signal output
rlabel metal3 s 519520 212984 520000 213104 6 gpio_dm1[10]
port 48 nsew signal output
rlabel metal3 s 519520 232568 520000 232688 6 gpio_dm1[11]
port 49 nsew signal output
rlabel metal3 s 519520 252152 520000 252272 6 gpio_dm1[12]
port 50 nsew signal output
rlabel metal3 s 519520 271736 520000 271856 6 gpio_dm1[13]
port 51 nsew signal output
rlabel metal3 s 519520 291320 520000 291440 6 gpio_dm1[14]
port 52 nsew signal output
rlabel metal2 s 506294 319520 506350 320000 6 gpio_dm1[15]
port 53 nsew signal output
rlabel metal2 s 448886 319520 448942 320000 6 gpio_dm1[16]
port 54 nsew signal output
rlabel metal2 s 391478 319520 391534 320000 6 gpio_dm1[17]
port 55 nsew signal output
rlabel metal2 s 334070 319520 334126 320000 6 gpio_dm1[18]
port 56 nsew signal output
rlabel metal2 s 276662 319520 276718 320000 6 gpio_dm1[19]
port 57 nsew signal output
rlabel metal3 s 519520 36728 520000 36848 6 gpio_dm1[1]
port 58 nsew signal output
rlabel metal2 s 219254 319520 219310 320000 6 gpio_dm1[20]
port 59 nsew signal output
rlabel metal2 s 161846 319520 161902 320000 6 gpio_dm1[21]
port 60 nsew signal output
rlabel metal2 s 104438 319520 104494 320000 6 gpio_dm1[22]
port 61 nsew signal output
rlabel metal2 s 47030 319520 47086 320000 6 gpio_dm1[23]
port 62 nsew signal output
rlabel metal3 s 0 294584 480 294704 6 gpio_dm1[24]
port 63 nsew signal output
rlabel metal3 s 0 275000 480 275120 6 gpio_dm1[25]
port 64 nsew signal output
rlabel metal3 s 0 255416 480 255536 6 gpio_dm1[26]
port 65 nsew signal output
rlabel metal3 s 0 235832 480 235952 6 gpio_dm1[27]
port 66 nsew signal output
rlabel metal3 s 0 216248 480 216368 6 gpio_dm1[28]
port 67 nsew signal output
rlabel metal3 s 0 196664 480 196784 6 gpio_dm1[29]
port 68 nsew signal output
rlabel metal3 s 519520 56312 520000 56432 6 gpio_dm1[2]
port 69 nsew signal output
rlabel metal3 s 0 177080 480 177200 6 gpio_dm1[30]
port 70 nsew signal output
rlabel metal3 s 0 157496 480 157616 6 gpio_dm1[31]
port 71 nsew signal output
rlabel metal3 s 0 137912 480 138032 6 gpio_dm1[32]
port 72 nsew signal output
rlabel metal3 s 0 118328 480 118448 6 gpio_dm1[33]
port 73 nsew signal output
rlabel metal3 s 0 98744 480 98864 6 gpio_dm1[34]
port 74 nsew signal output
rlabel metal3 s 0 79160 480 79280 6 gpio_dm1[35]
port 75 nsew signal output
rlabel metal3 s 0 59576 480 59696 6 gpio_dm1[36]
port 76 nsew signal output
rlabel metal3 s 0 39992 480 40112 6 gpio_dm1[37]
port 77 nsew signal output
rlabel metal2 s 20994 0 21050 480 6 gpio_dm1[38]
port 78 nsew signal output
rlabel metal2 s 79506 0 79562 480 6 gpio_dm1[39]
port 79 nsew signal output
rlabel metal3 s 519520 75896 520000 76016 6 gpio_dm1[3]
port 80 nsew signal output
rlabel metal2 s 138018 0 138074 480 6 gpio_dm1[40]
port 81 nsew signal output
rlabel metal2 s 196530 0 196586 480 6 gpio_dm1[41]
port 82 nsew signal output
rlabel metal2 s 255042 0 255098 480 6 gpio_dm1[42]
port 83 nsew signal output
rlabel metal2 s 313554 0 313610 480 6 gpio_dm1[43]
port 84 nsew signal output
rlabel metal3 s 519520 95480 520000 95600 6 gpio_dm1[4]
port 85 nsew signal output
rlabel metal3 s 519520 115064 520000 115184 6 gpio_dm1[5]
port 86 nsew signal output
rlabel metal3 s 519520 134648 520000 134768 6 gpio_dm1[6]
port 87 nsew signal output
rlabel metal3 s 519520 154232 520000 154352 6 gpio_dm1[7]
port 88 nsew signal output
rlabel metal3 s 519520 173816 520000 173936 6 gpio_dm1[8]
port 89 nsew signal output
rlabel metal3 s 519520 193400 520000 193520 6 gpio_dm1[9]
port 90 nsew signal output
rlabel metal3 s 519520 22040 520000 22160 6 gpio_dm2[0]
port 91 nsew signal output
rlabel metal3 s 519520 217880 520000 218000 6 gpio_dm2[10]
port 92 nsew signal output
rlabel metal3 s 519520 237464 520000 237584 6 gpio_dm2[11]
port 93 nsew signal output
rlabel metal3 s 519520 257048 520000 257168 6 gpio_dm2[12]
port 94 nsew signal output
rlabel metal3 s 519520 276632 520000 276752 6 gpio_dm2[13]
port 95 nsew signal output
rlabel metal3 s 519520 296216 520000 296336 6 gpio_dm2[14]
port 96 nsew signal output
rlabel metal2 s 491942 319520 491998 320000 6 gpio_dm2[15]
port 97 nsew signal output
rlabel metal2 s 434534 319520 434590 320000 6 gpio_dm2[16]
port 98 nsew signal output
rlabel metal2 s 377126 319520 377182 320000 6 gpio_dm2[17]
port 99 nsew signal output
rlabel metal2 s 319718 319520 319774 320000 6 gpio_dm2[18]
port 100 nsew signal output
rlabel metal2 s 262310 319520 262366 320000 6 gpio_dm2[19]
port 101 nsew signal output
rlabel metal3 s 519520 41624 520000 41744 6 gpio_dm2[1]
port 102 nsew signal output
rlabel metal2 s 204902 319520 204958 320000 6 gpio_dm2[20]
port 103 nsew signal output
rlabel metal2 s 147494 319520 147550 320000 6 gpio_dm2[21]
port 104 nsew signal output
rlabel metal2 s 90086 319520 90142 320000 6 gpio_dm2[22]
port 105 nsew signal output
rlabel metal2 s 32678 319520 32734 320000 6 gpio_dm2[23]
port 106 nsew signal output
rlabel metal3 s 0 289688 480 289808 6 gpio_dm2[24]
port 107 nsew signal output
rlabel metal3 s 0 270104 480 270224 6 gpio_dm2[25]
port 108 nsew signal output
rlabel metal3 s 0 250520 480 250640 6 gpio_dm2[26]
port 109 nsew signal output
rlabel metal3 s 0 230936 480 231056 6 gpio_dm2[27]
port 110 nsew signal output
rlabel metal3 s 0 211352 480 211472 6 gpio_dm2[28]
port 111 nsew signal output
rlabel metal3 s 0 191768 480 191888 6 gpio_dm2[29]
port 112 nsew signal output
rlabel metal3 s 519520 61208 520000 61328 6 gpio_dm2[2]
port 113 nsew signal output
rlabel metal3 s 0 172184 480 172304 6 gpio_dm2[30]
port 114 nsew signal output
rlabel metal3 s 0 152600 480 152720 6 gpio_dm2[31]
port 115 nsew signal output
rlabel metal3 s 0 133016 480 133136 6 gpio_dm2[32]
port 116 nsew signal output
rlabel metal3 s 0 113432 480 113552 6 gpio_dm2[33]
port 117 nsew signal output
rlabel metal3 s 0 93848 480 93968 6 gpio_dm2[34]
port 118 nsew signal output
rlabel metal3 s 0 74264 480 74384 6 gpio_dm2[35]
port 119 nsew signal output
rlabel metal3 s 0 54680 480 54800 6 gpio_dm2[36]
port 120 nsew signal output
rlabel metal3 s 0 35096 480 35216 6 gpio_dm2[37]
port 121 nsew signal output
rlabel metal2 s 35622 0 35678 480 6 gpio_dm2[38]
port 122 nsew signal output
rlabel metal2 s 94134 0 94190 480 6 gpio_dm2[39]
port 123 nsew signal output
rlabel metal3 s 519520 80792 520000 80912 6 gpio_dm2[3]
port 124 nsew signal output
rlabel metal2 s 152646 0 152702 480 6 gpio_dm2[40]
port 125 nsew signal output
rlabel metal2 s 211158 0 211214 480 6 gpio_dm2[41]
port 126 nsew signal output
rlabel metal2 s 269670 0 269726 480 6 gpio_dm2[42]
port 127 nsew signal output
rlabel metal2 s 328182 0 328238 480 6 gpio_dm2[43]
port 128 nsew signal output
rlabel metal3 s 519520 100376 520000 100496 6 gpio_dm2[4]
port 129 nsew signal output
rlabel metal3 s 519520 119960 520000 120080 6 gpio_dm2[5]
port 130 nsew signal output
rlabel metal3 s 519520 139544 520000 139664 6 gpio_dm2[6]
port 131 nsew signal output
rlabel metal3 s 519520 159128 520000 159248 6 gpio_dm2[7]
port 132 nsew signal output
rlabel metal3 s 519520 178712 520000 178832 6 gpio_dm2[8]
port 133 nsew signal output
rlabel metal3 s 519520 198296 520000 198416 6 gpio_dm2[9]
port 134 nsew signal output
rlabel metal3 s 519520 26936 520000 27056 6 gpio_ib_mode_sel[0]
port 135 nsew signal output
rlabel metal3 s 519520 222776 520000 222896 6 gpio_ib_mode_sel[10]
port 136 nsew signal output
rlabel metal3 s 519520 242360 520000 242480 6 gpio_ib_mode_sel[11]
port 137 nsew signal output
rlabel metal3 s 519520 261944 520000 262064 6 gpio_ib_mode_sel[12]
port 138 nsew signal output
rlabel metal3 s 519520 281528 520000 281648 6 gpio_ib_mode_sel[13]
port 139 nsew signal output
rlabel metal3 s 519520 301112 520000 301232 6 gpio_ib_mode_sel[14]
port 140 nsew signal output
rlabel metal2 s 477590 319520 477646 320000 6 gpio_ib_mode_sel[15]
port 141 nsew signal output
rlabel metal2 s 420182 319520 420238 320000 6 gpio_ib_mode_sel[16]
port 142 nsew signal output
rlabel metal2 s 362774 319520 362830 320000 6 gpio_ib_mode_sel[17]
port 143 nsew signal output
rlabel metal2 s 305366 319520 305422 320000 6 gpio_ib_mode_sel[18]
port 144 nsew signal output
rlabel metal2 s 247958 319520 248014 320000 6 gpio_ib_mode_sel[19]
port 145 nsew signal output
rlabel metal3 s 519520 46520 520000 46640 6 gpio_ib_mode_sel[1]
port 146 nsew signal output
rlabel metal2 s 190550 319520 190606 320000 6 gpio_ib_mode_sel[20]
port 147 nsew signal output
rlabel metal2 s 133142 319520 133198 320000 6 gpio_ib_mode_sel[21]
port 148 nsew signal output
rlabel metal2 s 75734 319520 75790 320000 6 gpio_ib_mode_sel[22]
port 149 nsew signal output
rlabel metal2 s 18326 319520 18382 320000 6 gpio_ib_mode_sel[23]
port 150 nsew signal output
rlabel metal3 s 0 284792 480 284912 6 gpio_ib_mode_sel[24]
port 151 nsew signal output
rlabel metal3 s 0 265208 480 265328 6 gpio_ib_mode_sel[25]
port 152 nsew signal output
rlabel metal3 s 0 245624 480 245744 6 gpio_ib_mode_sel[26]
port 153 nsew signal output
rlabel metal3 s 0 226040 480 226160 6 gpio_ib_mode_sel[27]
port 154 nsew signal output
rlabel metal3 s 0 206456 480 206576 6 gpio_ib_mode_sel[28]
port 155 nsew signal output
rlabel metal3 s 0 186872 480 186992 6 gpio_ib_mode_sel[29]
port 156 nsew signal output
rlabel metal3 s 519520 66104 520000 66224 6 gpio_ib_mode_sel[2]
port 157 nsew signal output
rlabel metal3 s 0 167288 480 167408 6 gpio_ib_mode_sel[30]
port 158 nsew signal output
rlabel metal3 s 0 147704 480 147824 6 gpio_ib_mode_sel[31]
port 159 nsew signal output
rlabel metal3 s 0 128120 480 128240 6 gpio_ib_mode_sel[32]
port 160 nsew signal output
rlabel metal3 s 0 108536 480 108656 6 gpio_ib_mode_sel[33]
port 161 nsew signal output
rlabel metal3 s 0 88952 480 89072 6 gpio_ib_mode_sel[34]
port 162 nsew signal output
rlabel metal3 s 0 69368 480 69488 6 gpio_ib_mode_sel[35]
port 163 nsew signal output
rlabel metal3 s 0 49784 480 49904 6 gpio_ib_mode_sel[36]
port 164 nsew signal output
rlabel metal3 s 0 30200 480 30320 6 gpio_ib_mode_sel[37]
port 165 nsew signal output
rlabel metal2 s 50250 0 50306 480 6 gpio_ib_mode_sel[38]
port 166 nsew signal output
rlabel metal2 s 108762 0 108818 480 6 gpio_ib_mode_sel[39]
port 167 nsew signal output
rlabel metal3 s 519520 85688 520000 85808 6 gpio_ib_mode_sel[3]
port 168 nsew signal output
rlabel metal2 s 167274 0 167330 480 6 gpio_ib_mode_sel[40]
port 169 nsew signal output
rlabel metal2 s 225786 0 225842 480 6 gpio_ib_mode_sel[41]
port 170 nsew signal output
rlabel metal2 s 284298 0 284354 480 6 gpio_ib_mode_sel[42]
port 171 nsew signal output
rlabel metal2 s 342810 0 342866 480 6 gpio_ib_mode_sel[43]
port 172 nsew signal output
rlabel metal3 s 519520 105272 520000 105392 6 gpio_ib_mode_sel[4]
port 173 nsew signal output
rlabel metal3 s 519520 124856 520000 124976 6 gpio_ib_mode_sel[5]
port 174 nsew signal output
rlabel metal3 s 519520 144440 520000 144560 6 gpio_ib_mode_sel[6]
port 175 nsew signal output
rlabel metal3 s 519520 164024 520000 164144 6 gpio_ib_mode_sel[7]
port 176 nsew signal output
rlabel metal3 s 519520 183608 520000 183728 6 gpio_ib_mode_sel[8]
port 177 nsew signal output
rlabel metal3 s 519520 203192 520000 203312 6 gpio_ib_mode_sel[9]
port 178 nsew signal output
rlabel metal3 s 519520 20408 520000 20528 6 gpio_ieb[0]
port 179 nsew signal output
rlabel metal3 s 519520 216248 520000 216368 6 gpio_ieb[10]
port 180 nsew signal output
rlabel metal3 s 519520 235832 520000 235952 6 gpio_ieb[11]
port 181 nsew signal output
rlabel metal3 s 519520 255416 520000 255536 6 gpio_ieb[12]
port 182 nsew signal output
rlabel metal3 s 519520 275000 520000 275120 6 gpio_ieb[13]
port 183 nsew signal output
rlabel metal3 s 519520 294584 520000 294704 6 gpio_ieb[14]
port 184 nsew signal output
rlabel metal2 s 496726 319520 496782 320000 6 gpio_ieb[15]
port 185 nsew signal output
rlabel metal2 s 439318 319520 439374 320000 6 gpio_ieb[16]
port 186 nsew signal output
rlabel metal2 s 381910 319520 381966 320000 6 gpio_ieb[17]
port 187 nsew signal output
rlabel metal2 s 324502 319520 324558 320000 6 gpio_ieb[18]
port 188 nsew signal output
rlabel metal2 s 267094 319520 267150 320000 6 gpio_ieb[19]
port 189 nsew signal output
rlabel metal3 s 519520 39992 520000 40112 6 gpio_ieb[1]
port 190 nsew signal output
rlabel metal2 s 209686 319520 209742 320000 6 gpio_ieb[20]
port 191 nsew signal output
rlabel metal2 s 152278 319520 152334 320000 6 gpio_ieb[21]
port 192 nsew signal output
rlabel metal2 s 94870 319520 94926 320000 6 gpio_ieb[22]
port 193 nsew signal output
rlabel metal2 s 37462 319520 37518 320000 6 gpio_ieb[23]
port 194 nsew signal output
rlabel metal3 s 0 291320 480 291440 6 gpio_ieb[24]
port 195 nsew signal output
rlabel metal3 s 0 271736 480 271856 6 gpio_ieb[25]
port 196 nsew signal output
rlabel metal3 s 0 252152 480 252272 6 gpio_ieb[26]
port 197 nsew signal output
rlabel metal3 s 0 232568 480 232688 6 gpio_ieb[27]
port 198 nsew signal output
rlabel metal3 s 0 212984 480 213104 6 gpio_ieb[28]
port 199 nsew signal output
rlabel metal3 s 0 193400 480 193520 6 gpio_ieb[29]
port 200 nsew signal output
rlabel metal3 s 519520 59576 520000 59696 6 gpio_ieb[2]
port 201 nsew signal output
rlabel metal3 s 0 173816 480 173936 6 gpio_ieb[30]
port 202 nsew signal output
rlabel metal3 s 0 154232 480 154352 6 gpio_ieb[31]
port 203 nsew signal output
rlabel metal3 s 0 134648 480 134768 6 gpio_ieb[32]
port 204 nsew signal output
rlabel metal3 s 0 115064 480 115184 6 gpio_ieb[33]
port 205 nsew signal output
rlabel metal3 s 0 95480 480 95600 6 gpio_ieb[34]
port 206 nsew signal output
rlabel metal3 s 0 75896 480 76016 6 gpio_ieb[35]
port 207 nsew signal output
rlabel metal3 s 0 56312 480 56432 6 gpio_ieb[36]
port 208 nsew signal output
rlabel metal3 s 0 36728 480 36848 6 gpio_ieb[37]
port 209 nsew signal output
rlabel metal2 s 30746 0 30802 480 6 gpio_ieb[38]
port 210 nsew signal output
rlabel metal2 s 89258 0 89314 480 6 gpio_ieb[39]
port 211 nsew signal output
rlabel metal3 s 519520 79160 520000 79280 6 gpio_ieb[3]
port 212 nsew signal output
rlabel metal2 s 147770 0 147826 480 6 gpio_ieb[40]
port 213 nsew signal output
rlabel metal2 s 206282 0 206338 480 6 gpio_ieb[41]
port 214 nsew signal output
rlabel metal2 s 264794 0 264850 480 6 gpio_ieb[42]
port 215 nsew signal output
rlabel metal2 s 323306 0 323362 480 6 gpio_ieb[43]
port 216 nsew signal output
rlabel metal3 s 519520 98744 520000 98864 6 gpio_ieb[4]
port 217 nsew signal output
rlabel metal3 s 519520 118328 520000 118448 6 gpio_ieb[5]
port 218 nsew signal output
rlabel metal3 s 519520 137912 520000 138032 6 gpio_ieb[6]
port 219 nsew signal output
rlabel metal3 s 519520 157496 520000 157616 6 gpio_ieb[7]
port 220 nsew signal output
rlabel metal3 s 519520 177080 520000 177200 6 gpio_ieb[8]
port 221 nsew signal output
rlabel metal3 s 519520 196664 520000 196784 6 gpio_ieb[9]
port 222 nsew signal output
rlabel metal3 s 519520 13880 520000 14000 6 gpio_in[0]
port 223 nsew signal input
rlabel metal3 s 519520 209720 520000 209840 6 gpio_in[10]
port 224 nsew signal input
rlabel metal3 s 519520 229304 520000 229424 6 gpio_in[11]
port 225 nsew signal input
rlabel metal3 s 519520 248888 520000 249008 6 gpio_in[12]
port 226 nsew signal input
rlabel metal3 s 519520 268472 520000 268592 6 gpio_in[13]
port 227 nsew signal input
rlabel metal3 s 519520 288056 520000 288176 6 gpio_in[14]
port 228 nsew signal input
rlabel metal2 s 515862 319520 515918 320000 6 gpio_in[15]
port 229 nsew signal input
rlabel metal2 s 458454 319520 458510 320000 6 gpio_in[16]
port 230 nsew signal input
rlabel metal2 s 401046 319520 401102 320000 6 gpio_in[17]
port 231 nsew signal input
rlabel metal2 s 343638 319520 343694 320000 6 gpio_in[18]
port 232 nsew signal input
rlabel metal2 s 286230 319520 286286 320000 6 gpio_in[19]
port 233 nsew signal input
rlabel metal3 s 519520 33464 520000 33584 6 gpio_in[1]
port 234 nsew signal input
rlabel metal2 s 228822 319520 228878 320000 6 gpio_in[20]
port 235 nsew signal input
rlabel metal2 s 171414 319520 171470 320000 6 gpio_in[21]
port 236 nsew signal input
rlabel metal2 s 114006 319520 114062 320000 6 gpio_in[22]
port 237 nsew signal input
rlabel metal2 s 56598 319520 56654 320000 6 gpio_in[23]
port 238 nsew signal input
rlabel metal3 s 0 297848 480 297968 6 gpio_in[24]
port 239 nsew signal input
rlabel metal3 s 0 278264 480 278384 6 gpio_in[25]
port 240 nsew signal input
rlabel metal3 s 0 258680 480 258800 6 gpio_in[26]
port 241 nsew signal input
rlabel metal3 s 0 239096 480 239216 6 gpio_in[27]
port 242 nsew signal input
rlabel metal3 s 0 219512 480 219632 6 gpio_in[28]
port 243 nsew signal input
rlabel metal3 s 0 199928 480 200048 6 gpio_in[29]
port 244 nsew signal input
rlabel metal3 s 519520 53048 520000 53168 6 gpio_in[2]
port 245 nsew signal input
rlabel metal3 s 0 180344 480 180464 6 gpio_in[30]
port 246 nsew signal input
rlabel metal3 s 0 160760 480 160880 6 gpio_in[31]
port 247 nsew signal input
rlabel metal3 s 0 141176 480 141296 6 gpio_in[32]
port 248 nsew signal input
rlabel metal3 s 0 121592 480 121712 6 gpio_in[33]
port 249 nsew signal input
rlabel metal3 s 0 102008 480 102128 6 gpio_in[34]
port 250 nsew signal input
rlabel metal3 s 0 82424 480 82544 6 gpio_in[35]
port 251 nsew signal input
rlabel metal3 s 0 62840 480 62960 6 gpio_in[36]
port 252 nsew signal input
rlabel metal3 s 0 43256 480 43376 6 gpio_in[37]
port 253 nsew signal input
rlabel metal2 s 11242 0 11298 480 6 gpio_in[38]
port 254 nsew signal input
rlabel metal2 s 69754 0 69810 480 6 gpio_in[39]
port 255 nsew signal input
rlabel metal3 s 519520 72632 520000 72752 6 gpio_in[3]
port 256 nsew signal input
rlabel metal2 s 128266 0 128322 480 6 gpio_in[40]
port 257 nsew signal input
rlabel metal2 s 186778 0 186834 480 6 gpio_in[41]
port 258 nsew signal input
rlabel metal2 s 245290 0 245346 480 6 gpio_in[42]
port 259 nsew signal input
rlabel metal2 s 303802 0 303858 480 6 gpio_in[43]
port 260 nsew signal input
rlabel metal3 s 519520 92216 520000 92336 6 gpio_in[4]
port 261 nsew signal input
rlabel metal3 s 519520 111800 520000 111920 6 gpio_in[5]
port 262 nsew signal input
rlabel metal3 s 519520 131384 520000 131504 6 gpio_in[6]
port 263 nsew signal input
rlabel metal3 s 519520 150968 520000 151088 6 gpio_in[7]
port 264 nsew signal input
rlabel metal3 s 519520 170552 520000 170672 6 gpio_in[8]
port 265 nsew signal input
rlabel metal3 s 519520 190136 520000 190256 6 gpio_in[9]
port 266 nsew signal input
rlabel metal3 s 519520 30200 520000 30320 6 gpio_loopback_one[0]
port 267 nsew signal input
rlabel metal3 s 519520 226040 520000 226160 6 gpio_loopback_one[10]
port 268 nsew signal input
rlabel metal3 s 519520 245624 520000 245744 6 gpio_loopback_one[11]
port 269 nsew signal input
rlabel metal3 s 519520 265208 520000 265328 6 gpio_loopback_one[12]
port 270 nsew signal input
rlabel metal3 s 519520 284792 520000 284912 6 gpio_loopback_one[13]
port 271 nsew signal input
rlabel metal3 s 519520 304376 520000 304496 6 gpio_loopback_one[14]
port 272 nsew signal input
rlabel metal2 s 468022 319520 468078 320000 6 gpio_loopback_one[15]
port 273 nsew signal input
rlabel metal2 s 410614 319520 410670 320000 6 gpio_loopback_one[16]
port 274 nsew signal input
rlabel metal2 s 353206 319520 353262 320000 6 gpio_loopback_one[17]
port 275 nsew signal input
rlabel metal2 s 295798 319520 295854 320000 6 gpio_loopback_one[18]
port 276 nsew signal input
rlabel metal2 s 238390 319520 238446 320000 6 gpio_loopback_one[19]
port 277 nsew signal input
rlabel metal3 s 519520 49784 520000 49904 6 gpio_loopback_one[1]
port 278 nsew signal input
rlabel metal2 s 180982 319520 181038 320000 6 gpio_loopback_one[20]
port 279 nsew signal input
rlabel metal2 s 123574 319520 123630 320000 6 gpio_loopback_one[21]
port 280 nsew signal input
rlabel metal2 s 66166 319520 66222 320000 6 gpio_loopback_one[22]
port 281 nsew signal input
rlabel metal2 s 8758 319520 8814 320000 6 gpio_loopback_one[23]
port 282 nsew signal input
rlabel metal3 s 0 281528 480 281648 6 gpio_loopback_one[24]
port 283 nsew signal input
rlabel metal3 s 0 261944 480 262064 6 gpio_loopback_one[25]
port 284 nsew signal input
rlabel metal3 s 0 242360 480 242480 6 gpio_loopback_one[26]
port 285 nsew signal input
rlabel metal3 s 0 222776 480 222896 6 gpio_loopback_one[27]
port 286 nsew signal input
rlabel metal3 s 0 203192 480 203312 6 gpio_loopback_one[28]
port 287 nsew signal input
rlabel metal3 s 0 183608 480 183728 6 gpio_loopback_one[29]
port 288 nsew signal input
rlabel metal3 s 519520 69368 520000 69488 6 gpio_loopback_one[2]
port 289 nsew signal input
rlabel metal3 s 0 164024 480 164144 6 gpio_loopback_one[30]
port 290 nsew signal input
rlabel metal3 s 0 144440 480 144560 6 gpio_loopback_one[31]
port 291 nsew signal input
rlabel metal3 s 0 124856 480 124976 6 gpio_loopback_one[32]
port 292 nsew signal input
rlabel metal3 s 0 105272 480 105392 6 gpio_loopback_one[33]
port 293 nsew signal input
rlabel metal3 s 0 85688 480 85808 6 gpio_loopback_one[34]
port 294 nsew signal input
rlabel metal3 s 0 66104 480 66224 6 gpio_loopback_one[35]
port 295 nsew signal input
rlabel metal3 s 0 46520 480 46640 6 gpio_loopback_one[36]
port 296 nsew signal input
rlabel metal3 s 0 26936 480 27056 6 gpio_loopback_one[37]
port 297 nsew signal input
rlabel metal2 s 60002 0 60058 480 6 gpio_loopback_one[38]
port 298 nsew signal input
rlabel metal2 s 118514 0 118570 480 6 gpio_loopback_one[39]
port 299 nsew signal input
rlabel metal3 s 519520 88952 520000 89072 6 gpio_loopback_one[3]
port 300 nsew signal input
rlabel metal2 s 177026 0 177082 480 6 gpio_loopback_one[40]
port 301 nsew signal input
rlabel metal2 s 235538 0 235594 480 6 gpio_loopback_one[41]
port 302 nsew signal input
rlabel metal2 s 294050 0 294106 480 6 gpio_loopback_one[42]
port 303 nsew signal input
rlabel metal2 s 352562 0 352618 480 6 gpio_loopback_one[43]
port 304 nsew signal input
rlabel metal3 s 519520 108536 520000 108656 6 gpio_loopback_one[4]
port 305 nsew signal input
rlabel metal3 s 519520 128120 520000 128240 6 gpio_loopback_one[5]
port 306 nsew signal input
rlabel metal3 s 519520 147704 520000 147824 6 gpio_loopback_one[6]
port 307 nsew signal input
rlabel metal3 s 519520 167288 520000 167408 6 gpio_loopback_one[7]
port 308 nsew signal input
rlabel metal3 s 519520 186872 520000 186992 6 gpio_loopback_one[8]
port 309 nsew signal input
rlabel metal3 s 519520 206456 520000 206576 6 gpio_loopback_one[9]
port 310 nsew signal input
rlabel metal3 s 519520 31832 520000 31952 6 gpio_loopback_zero[0]
port 311 nsew signal input
rlabel metal3 s 519520 227672 520000 227792 6 gpio_loopback_zero[10]
port 312 nsew signal input
rlabel metal3 s 519520 247256 520000 247376 6 gpio_loopback_zero[11]
port 313 nsew signal input
rlabel metal3 s 519520 266840 520000 266960 6 gpio_loopback_zero[12]
port 314 nsew signal input
rlabel metal3 s 519520 286424 520000 286544 6 gpio_loopback_zero[13]
port 315 nsew signal input
rlabel metal3 s 519520 306008 520000 306128 6 gpio_loopback_zero[14]
port 316 nsew signal input
rlabel metal2 s 463238 319520 463294 320000 6 gpio_loopback_zero[15]
port 317 nsew signal input
rlabel metal2 s 405830 319520 405886 320000 6 gpio_loopback_zero[16]
port 318 nsew signal input
rlabel metal2 s 348422 319520 348478 320000 6 gpio_loopback_zero[17]
port 319 nsew signal input
rlabel metal2 s 291014 319520 291070 320000 6 gpio_loopback_zero[18]
port 320 nsew signal input
rlabel metal2 s 233606 319520 233662 320000 6 gpio_loopback_zero[19]
port 321 nsew signal input
rlabel metal3 s 519520 51416 520000 51536 6 gpio_loopback_zero[1]
port 322 nsew signal input
rlabel metal2 s 176198 319520 176254 320000 6 gpio_loopback_zero[20]
port 323 nsew signal input
rlabel metal2 s 118790 319520 118846 320000 6 gpio_loopback_zero[21]
port 324 nsew signal input
rlabel metal2 s 61382 319520 61438 320000 6 gpio_loopback_zero[22]
port 325 nsew signal input
rlabel metal2 s 3974 319520 4030 320000 6 gpio_loopback_zero[23]
port 326 nsew signal input
rlabel metal3 s 0 279896 480 280016 6 gpio_loopback_zero[24]
port 327 nsew signal input
rlabel metal3 s 0 260312 480 260432 6 gpio_loopback_zero[25]
port 328 nsew signal input
rlabel metal3 s 0 240728 480 240848 6 gpio_loopback_zero[26]
port 329 nsew signal input
rlabel metal3 s 0 221144 480 221264 6 gpio_loopback_zero[27]
port 330 nsew signal input
rlabel metal3 s 0 201560 480 201680 6 gpio_loopback_zero[28]
port 331 nsew signal input
rlabel metal3 s 0 181976 480 182096 6 gpio_loopback_zero[29]
port 332 nsew signal input
rlabel metal3 s 519520 71000 520000 71120 6 gpio_loopback_zero[2]
port 333 nsew signal input
rlabel metal3 s 0 162392 480 162512 6 gpio_loopback_zero[30]
port 334 nsew signal input
rlabel metal3 s 0 142808 480 142928 6 gpio_loopback_zero[31]
port 335 nsew signal input
rlabel metal3 s 0 123224 480 123344 6 gpio_loopback_zero[32]
port 336 nsew signal input
rlabel metal3 s 0 103640 480 103760 6 gpio_loopback_zero[33]
port 337 nsew signal input
rlabel metal3 s 0 84056 480 84176 6 gpio_loopback_zero[34]
port 338 nsew signal input
rlabel metal3 s 0 64472 480 64592 6 gpio_loopback_zero[35]
port 339 nsew signal input
rlabel metal3 s 0 44888 480 45008 6 gpio_loopback_zero[36]
port 340 nsew signal input
rlabel metal3 s 0 25304 480 25424 6 gpio_loopback_zero[37]
port 341 nsew signal input
rlabel metal2 s 64878 0 64934 480 6 gpio_loopback_zero[38]
port 342 nsew signal input
rlabel metal2 s 123390 0 123446 480 6 gpio_loopback_zero[39]
port 343 nsew signal input
rlabel metal3 s 519520 90584 520000 90704 6 gpio_loopback_zero[3]
port 344 nsew signal input
rlabel metal2 s 181902 0 181958 480 6 gpio_loopback_zero[40]
port 345 nsew signal input
rlabel metal2 s 240414 0 240470 480 6 gpio_loopback_zero[41]
port 346 nsew signal input
rlabel metal2 s 298926 0 298982 480 6 gpio_loopback_zero[42]
port 347 nsew signal input
rlabel metal2 s 357438 0 357494 480 6 gpio_loopback_zero[43]
port 348 nsew signal input
rlabel metal3 s 519520 110168 520000 110288 6 gpio_loopback_zero[4]
port 349 nsew signal input
rlabel metal3 s 519520 129752 520000 129872 6 gpio_loopback_zero[5]
port 350 nsew signal input
rlabel metal3 s 519520 149336 520000 149456 6 gpio_loopback_zero[6]
port 351 nsew signal input
rlabel metal3 s 519520 168920 520000 169040 6 gpio_loopback_zero[7]
port 352 nsew signal input
rlabel metal3 s 519520 188504 520000 188624 6 gpio_loopback_zero[8]
port 353 nsew signal input
rlabel metal3 s 519520 208088 520000 208208 6 gpio_loopback_zero[9]
port 354 nsew signal input
rlabel metal3 s 519520 28568 520000 28688 6 gpio_oeb[0]
port 355 nsew signal output
rlabel metal3 s 519520 224408 520000 224528 6 gpio_oeb[10]
port 356 nsew signal output
rlabel metal3 s 519520 243992 520000 244112 6 gpio_oeb[11]
port 357 nsew signal output
rlabel metal3 s 519520 263576 520000 263696 6 gpio_oeb[12]
port 358 nsew signal output
rlabel metal3 s 519520 283160 520000 283280 6 gpio_oeb[13]
port 359 nsew signal output
rlabel metal3 s 519520 302744 520000 302864 6 gpio_oeb[14]
port 360 nsew signal output
rlabel metal2 s 472806 319520 472862 320000 6 gpio_oeb[15]
port 361 nsew signal output
rlabel metal2 s 415398 319520 415454 320000 6 gpio_oeb[16]
port 362 nsew signal output
rlabel metal2 s 357990 319520 358046 320000 6 gpio_oeb[17]
port 363 nsew signal output
rlabel metal2 s 300582 319520 300638 320000 6 gpio_oeb[18]
port 364 nsew signal output
rlabel metal2 s 243174 319520 243230 320000 6 gpio_oeb[19]
port 365 nsew signal output
rlabel metal3 s 519520 48152 520000 48272 6 gpio_oeb[1]
port 366 nsew signal output
rlabel metal2 s 185766 319520 185822 320000 6 gpio_oeb[20]
port 367 nsew signal output
rlabel metal2 s 128358 319520 128414 320000 6 gpio_oeb[21]
port 368 nsew signal output
rlabel metal2 s 70950 319520 71006 320000 6 gpio_oeb[22]
port 369 nsew signal output
rlabel metal2 s 13542 319520 13598 320000 6 gpio_oeb[23]
port 370 nsew signal output
rlabel metal3 s 0 283160 480 283280 6 gpio_oeb[24]
port 371 nsew signal output
rlabel metal3 s 0 263576 480 263696 6 gpio_oeb[25]
port 372 nsew signal output
rlabel metal3 s 0 243992 480 244112 6 gpio_oeb[26]
port 373 nsew signal output
rlabel metal3 s 0 224408 480 224528 6 gpio_oeb[27]
port 374 nsew signal output
rlabel metal3 s 0 204824 480 204944 6 gpio_oeb[28]
port 375 nsew signal output
rlabel metal3 s 0 185240 480 185360 6 gpio_oeb[29]
port 376 nsew signal output
rlabel metal3 s 519520 67736 520000 67856 6 gpio_oeb[2]
port 377 nsew signal output
rlabel metal3 s 0 165656 480 165776 6 gpio_oeb[30]
port 378 nsew signal output
rlabel metal3 s 0 146072 480 146192 6 gpio_oeb[31]
port 379 nsew signal output
rlabel metal3 s 0 126488 480 126608 6 gpio_oeb[32]
port 380 nsew signal output
rlabel metal3 s 0 106904 480 107024 6 gpio_oeb[33]
port 381 nsew signal output
rlabel metal3 s 0 87320 480 87440 6 gpio_oeb[34]
port 382 nsew signal output
rlabel metal3 s 0 67736 480 67856 6 gpio_oeb[35]
port 383 nsew signal output
rlabel metal3 s 0 48152 480 48272 6 gpio_oeb[36]
port 384 nsew signal output
rlabel metal3 s 0 28568 480 28688 6 gpio_oeb[37]
port 385 nsew signal output
rlabel metal2 s 55126 0 55182 480 6 gpio_oeb[38]
port 386 nsew signal output
rlabel metal2 s 113638 0 113694 480 6 gpio_oeb[39]
port 387 nsew signal output
rlabel metal3 s 519520 87320 520000 87440 6 gpio_oeb[3]
port 388 nsew signal output
rlabel metal2 s 172150 0 172206 480 6 gpio_oeb[40]
port 389 nsew signal output
rlabel metal2 s 230662 0 230718 480 6 gpio_oeb[41]
port 390 nsew signal output
rlabel metal2 s 289174 0 289230 480 6 gpio_oeb[42]
port 391 nsew signal output
rlabel metal2 s 347686 0 347742 480 6 gpio_oeb[43]
port 392 nsew signal output
rlabel metal3 s 519520 106904 520000 107024 6 gpio_oeb[4]
port 393 nsew signal output
rlabel metal3 s 519520 126488 520000 126608 6 gpio_oeb[5]
port 394 nsew signal output
rlabel metal3 s 519520 146072 520000 146192 6 gpio_oeb[6]
port 395 nsew signal output
rlabel metal3 s 519520 165656 520000 165776 6 gpio_oeb[7]
port 396 nsew signal output
rlabel metal3 s 519520 185240 520000 185360 6 gpio_oeb[8]
port 397 nsew signal output
rlabel metal3 s 519520 204824 520000 204944 6 gpio_oeb[9]
port 398 nsew signal output
rlabel metal3 s 519520 23672 520000 23792 6 gpio_out[0]
port 399 nsew signal output
rlabel metal3 s 519520 219512 520000 219632 6 gpio_out[10]
port 400 nsew signal output
rlabel metal3 s 519520 239096 520000 239216 6 gpio_out[11]
port 401 nsew signal output
rlabel metal3 s 519520 258680 520000 258800 6 gpio_out[12]
port 402 nsew signal output
rlabel metal3 s 519520 278264 520000 278384 6 gpio_out[13]
port 403 nsew signal output
rlabel metal3 s 519520 297848 520000 297968 6 gpio_out[14]
port 404 nsew signal output
rlabel metal2 s 487158 319520 487214 320000 6 gpio_out[15]
port 405 nsew signal output
rlabel metal2 s 429750 319520 429806 320000 6 gpio_out[16]
port 406 nsew signal output
rlabel metal2 s 372342 319520 372398 320000 6 gpio_out[17]
port 407 nsew signal output
rlabel metal2 s 314934 319520 314990 320000 6 gpio_out[18]
port 408 nsew signal output
rlabel metal2 s 257526 319520 257582 320000 6 gpio_out[19]
port 409 nsew signal output
rlabel metal3 s 519520 43256 520000 43376 6 gpio_out[1]
port 410 nsew signal output
rlabel metal2 s 200118 319520 200174 320000 6 gpio_out[20]
port 411 nsew signal output
rlabel metal2 s 142710 319520 142766 320000 6 gpio_out[21]
port 412 nsew signal output
rlabel metal2 s 85302 319520 85358 320000 6 gpio_out[22]
port 413 nsew signal output
rlabel metal2 s 27894 319520 27950 320000 6 gpio_out[23]
port 414 nsew signal output
rlabel metal3 s 0 288056 480 288176 6 gpio_out[24]
port 415 nsew signal output
rlabel metal3 s 0 268472 480 268592 6 gpio_out[25]
port 416 nsew signal output
rlabel metal3 s 0 248888 480 249008 6 gpio_out[26]
port 417 nsew signal output
rlabel metal3 s 0 229304 480 229424 6 gpio_out[27]
port 418 nsew signal output
rlabel metal3 s 0 209720 480 209840 6 gpio_out[28]
port 419 nsew signal output
rlabel metal3 s 0 190136 480 190256 6 gpio_out[29]
port 420 nsew signal output
rlabel metal3 s 519520 62840 520000 62960 6 gpio_out[2]
port 421 nsew signal output
rlabel metal3 s 0 170552 480 170672 6 gpio_out[30]
port 422 nsew signal output
rlabel metal3 s 0 150968 480 151088 6 gpio_out[31]
port 423 nsew signal output
rlabel metal3 s 0 131384 480 131504 6 gpio_out[32]
port 424 nsew signal output
rlabel metal3 s 0 111800 480 111920 6 gpio_out[33]
port 425 nsew signal output
rlabel metal3 s 0 92216 480 92336 6 gpio_out[34]
port 426 nsew signal output
rlabel metal3 s 0 72632 480 72752 6 gpio_out[35]
port 427 nsew signal output
rlabel metal3 s 0 53048 480 53168 6 gpio_out[36]
port 428 nsew signal output
rlabel metal3 s 0 33464 480 33584 6 gpio_out[37]
port 429 nsew signal output
rlabel metal2 s 40498 0 40554 480 6 gpio_out[38]
port 430 nsew signal output
rlabel metal2 s 99010 0 99066 480 6 gpio_out[39]
port 431 nsew signal output
rlabel metal3 s 519520 82424 520000 82544 6 gpio_out[3]
port 432 nsew signal output
rlabel metal2 s 157522 0 157578 480 6 gpio_out[40]
port 433 nsew signal output
rlabel metal2 s 216034 0 216090 480 6 gpio_out[41]
port 434 nsew signal output
rlabel metal2 s 274546 0 274602 480 6 gpio_out[42]
port 435 nsew signal output
rlabel metal2 s 333058 0 333114 480 6 gpio_out[43]
port 436 nsew signal output
rlabel metal3 s 519520 102008 520000 102128 6 gpio_out[4]
port 437 nsew signal output
rlabel metal3 s 519520 121592 520000 121712 6 gpio_out[5]
port 438 nsew signal output
rlabel metal3 s 519520 141176 520000 141296 6 gpio_out[6]
port 439 nsew signal output
rlabel metal3 s 519520 160760 520000 160880 6 gpio_out[7]
port 440 nsew signal output
rlabel metal3 s 519520 180344 520000 180464 6 gpio_out[8]
port 441 nsew signal output
rlabel metal3 s 519520 199928 520000 200048 6 gpio_out[9]
port 442 nsew signal output
rlabel metal3 s 519520 15512 520000 15632 6 gpio_slow_sel[0]
port 443 nsew signal output
rlabel metal3 s 519520 211352 520000 211472 6 gpio_slow_sel[10]
port 444 nsew signal output
rlabel metal3 s 519520 230936 520000 231056 6 gpio_slow_sel[11]
port 445 nsew signal output
rlabel metal3 s 519520 250520 520000 250640 6 gpio_slow_sel[12]
port 446 nsew signal output
rlabel metal3 s 519520 270104 520000 270224 6 gpio_slow_sel[13]
port 447 nsew signal output
rlabel metal3 s 519520 289688 520000 289808 6 gpio_slow_sel[14]
port 448 nsew signal output
rlabel metal2 s 511078 319520 511134 320000 6 gpio_slow_sel[15]
port 449 nsew signal output
rlabel metal2 s 453670 319520 453726 320000 6 gpio_slow_sel[16]
port 450 nsew signal output
rlabel metal2 s 396262 319520 396318 320000 6 gpio_slow_sel[17]
port 451 nsew signal output
rlabel metal2 s 338854 319520 338910 320000 6 gpio_slow_sel[18]
port 452 nsew signal output
rlabel metal2 s 281446 319520 281502 320000 6 gpio_slow_sel[19]
port 453 nsew signal output
rlabel metal3 s 519520 35096 520000 35216 6 gpio_slow_sel[1]
port 454 nsew signal output
rlabel metal2 s 224038 319520 224094 320000 6 gpio_slow_sel[20]
port 455 nsew signal output
rlabel metal2 s 166630 319520 166686 320000 6 gpio_slow_sel[21]
port 456 nsew signal output
rlabel metal2 s 109222 319520 109278 320000 6 gpio_slow_sel[22]
port 457 nsew signal output
rlabel metal2 s 51814 319520 51870 320000 6 gpio_slow_sel[23]
port 458 nsew signal output
rlabel metal3 s 0 296216 480 296336 6 gpio_slow_sel[24]
port 459 nsew signal output
rlabel metal3 s 0 276632 480 276752 6 gpio_slow_sel[25]
port 460 nsew signal output
rlabel metal3 s 0 257048 480 257168 6 gpio_slow_sel[26]
port 461 nsew signal output
rlabel metal3 s 0 237464 480 237584 6 gpio_slow_sel[27]
port 462 nsew signal output
rlabel metal3 s 0 217880 480 218000 6 gpio_slow_sel[28]
port 463 nsew signal output
rlabel metal3 s 0 198296 480 198416 6 gpio_slow_sel[29]
port 464 nsew signal output
rlabel metal3 s 519520 54680 520000 54800 6 gpio_slow_sel[2]
port 465 nsew signal output
rlabel metal3 s 0 178712 480 178832 6 gpio_slow_sel[30]
port 466 nsew signal output
rlabel metal3 s 0 159128 480 159248 6 gpio_slow_sel[31]
port 467 nsew signal output
rlabel metal3 s 0 139544 480 139664 6 gpio_slow_sel[32]
port 468 nsew signal output
rlabel metal3 s 0 119960 480 120080 6 gpio_slow_sel[33]
port 469 nsew signal output
rlabel metal3 s 0 100376 480 100496 6 gpio_slow_sel[34]
port 470 nsew signal output
rlabel metal3 s 0 80792 480 80912 6 gpio_slow_sel[35]
port 471 nsew signal output
rlabel metal3 s 0 61208 480 61328 6 gpio_slow_sel[36]
port 472 nsew signal output
rlabel metal3 s 0 41624 480 41744 6 gpio_slow_sel[37]
port 473 nsew signal output
rlabel metal2 s 16118 0 16174 480 6 gpio_slow_sel[38]
port 474 nsew signal output
rlabel metal2 s 74630 0 74686 480 6 gpio_slow_sel[39]
port 475 nsew signal output
rlabel metal3 s 519520 74264 520000 74384 6 gpio_slow_sel[3]
port 476 nsew signal output
rlabel metal2 s 133142 0 133198 480 6 gpio_slow_sel[40]
port 477 nsew signal output
rlabel metal2 s 191654 0 191710 480 6 gpio_slow_sel[41]
port 478 nsew signal output
rlabel metal2 s 250166 0 250222 480 6 gpio_slow_sel[42]
port 479 nsew signal output
rlabel metal2 s 308678 0 308734 480 6 gpio_slow_sel[43]
port 480 nsew signal output
rlabel metal3 s 519520 93848 520000 93968 6 gpio_slow_sel[4]
port 481 nsew signal output
rlabel metal3 s 519520 113432 520000 113552 6 gpio_slow_sel[5]
port 482 nsew signal output
rlabel metal3 s 519520 133016 520000 133136 6 gpio_slow_sel[6]
port 483 nsew signal output
rlabel metal3 s 519520 152600 520000 152720 6 gpio_slow_sel[7]
port 484 nsew signal output
rlabel metal3 s 519520 172184 520000 172304 6 gpio_slow_sel[8]
port 485 nsew signal output
rlabel metal3 s 519520 191768 520000 191888 6 gpio_slow_sel[9]
port 486 nsew signal output
rlabel metal3 s 519520 25304 520000 25424 6 gpio_vtrip_sel[0]
port 487 nsew signal output
rlabel metal3 s 519520 221144 520000 221264 6 gpio_vtrip_sel[10]
port 488 nsew signal output
rlabel metal3 s 519520 240728 520000 240848 6 gpio_vtrip_sel[11]
port 489 nsew signal output
rlabel metal3 s 519520 260312 520000 260432 6 gpio_vtrip_sel[12]
port 490 nsew signal output
rlabel metal3 s 519520 279896 520000 280016 6 gpio_vtrip_sel[13]
port 491 nsew signal output
rlabel metal3 s 519520 299480 520000 299600 6 gpio_vtrip_sel[14]
port 492 nsew signal output
rlabel metal2 s 482374 319520 482430 320000 6 gpio_vtrip_sel[15]
port 493 nsew signal output
rlabel metal2 s 424966 319520 425022 320000 6 gpio_vtrip_sel[16]
port 494 nsew signal output
rlabel metal2 s 367558 319520 367614 320000 6 gpio_vtrip_sel[17]
port 495 nsew signal output
rlabel metal2 s 310150 319520 310206 320000 6 gpio_vtrip_sel[18]
port 496 nsew signal output
rlabel metal2 s 252742 319520 252798 320000 6 gpio_vtrip_sel[19]
port 497 nsew signal output
rlabel metal3 s 519520 44888 520000 45008 6 gpio_vtrip_sel[1]
port 498 nsew signal output
rlabel metal2 s 195334 319520 195390 320000 6 gpio_vtrip_sel[20]
port 499 nsew signal output
rlabel metal2 s 137926 319520 137982 320000 6 gpio_vtrip_sel[21]
port 500 nsew signal output
rlabel metal2 s 80518 319520 80574 320000 6 gpio_vtrip_sel[22]
port 501 nsew signal output
rlabel metal2 s 23110 319520 23166 320000 6 gpio_vtrip_sel[23]
port 502 nsew signal output
rlabel metal3 s 0 286424 480 286544 6 gpio_vtrip_sel[24]
port 503 nsew signal output
rlabel metal3 s 0 266840 480 266960 6 gpio_vtrip_sel[25]
port 504 nsew signal output
rlabel metal3 s 0 247256 480 247376 6 gpio_vtrip_sel[26]
port 505 nsew signal output
rlabel metal3 s 0 227672 480 227792 6 gpio_vtrip_sel[27]
port 506 nsew signal output
rlabel metal3 s 0 208088 480 208208 6 gpio_vtrip_sel[28]
port 507 nsew signal output
rlabel metal3 s 0 188504 480 188624 6 gpio_vtrip_sel[29]
port 508 nsew signal output
rlabel metal3 s 519520 64472 520000 64592 6 gpio_vtrip_sel[2]
port 509 nsew signal output
rlabel metal3 s 0 168920 480 169040 6 gpio_vtrip_sel[30]
port 510 nsew signal output
rlabel metal3 s 0 149336 480 149456 6 gpio_vtrip_sel[31]
port 511 nsew signal output
rlabel metal3 s 0 129752 480 129872 6 gpio_vtrip_sel[32]
port 512 nsew signal output
rlabel metal3 s 0 110168 480 110288 6 gpio_vtrip_sel[33]
port 513 nsew signal output
rlabel metal3 s 0 90584 480 90704 6 gpio_vtrip_sel[34]
port 514 nsew signal output
rlabel metal3 s 0 71000 480 71120 6 gpio_vtrip_sel[35]
port 515 nsew signal output
rlabel metal3 s 0 51416 480 51536 6 gpio_vtrip_sel[36]
port 516 nsew signal output
rlabel metal3 s 0 31832 480 31952 6 gpio_vtrip_sel[37]
port 517 nsew signal output
rlabel metal2 s 45374 0 45430 480 6 gpio_vtrip_sel[38]
port 518 nsew signal output
rlabel metal2 s 103886 0 103942 480 6 gpio_vtrip_sel[39]
port 519 nsew signal output
rlabel metal3 s 519520 84056 520000 84176 6 gpio_vtrip_sel[3]
port 520 nsew signal output
rlabel metal2 s 162398 0 162454 480 6 gpio_vtrip_sel[40]
port 521 nsew signal output
rlabel metal2 s 220910 0 220966 480 6 gpio_vtrip_sel[41]
port 522 nsew signal output
rlabel metal2 s 279422 0 279478 480 6 gpio_vtrip_sel[42]
port 523 nsew signal output
rlabel metal2 s 337934 0 337990 480 6 gpio_vtrip_sel[43]
port 524 nsew signal output
rlabel metal3 s 519520 103640 520000 103760 6 gpio_vtrip_sel[4]
port 525 nsew signal output
rlabel metal3 s 519520 123224 520000 123344 6 gpio_vtrip_sel[5]
port 526 nsew signal output
rlabel metal3 s 519520 142808 520000 142928 6 gpio_vtrip_sel[6]
port 527 nsew signal output
rlabel metal3 s 519520 162392 520000 162512 6 gpio_vtrip_sel[7]
port 528 nsew signal output
rlabel metal3 s 519520 181976 520000 182096 6 gpio_vtrip_sel[8]
port 529 nsew signal output
rlabel metal3 s 519520 201560 520000 201680 6 gpio_vtrip_sel[9]
port 530 nsew signal output
rlabel metal2 s 362314 0 362370 480 6 mask_rev[0]
port 531 nsew signal input
rlabel metal2 s 411074 0 411130 480 6 mask_rev[10]
port 532 nsew signal input
rlabel metal2 s 415950 0 416006 480 6 mask_rev[11]
port 533 nsew signal input
rlabel metal2 s 420826 0 420882 480 6 mask_rev[12]
port 534 nsew signal input
rlabel metal2 s 425702 0 425758 480 6 mask_rev[13]
port 535 nsew signal input
rlabel metal2 s 430578 0 430634 480 6 mask_rev[14]
port 536 nsew signal input
rlabel metal2 s 435454 0 435510 480 6 mask_rev[15]
port 537 nsew signal input
rlabel metal2 s 440330 0 440386 480 6 mask_rev[16]
port 538 nsew signal input
rlabel metal2 s 445206 0 445262 480 6 mask_rev[17]
port 539 nsew signal input
rlabel metal2 s 450082 0 450138 480 6 mask_rev[18]
port 540 nsew signal input
rlabel metal2 s 454958 0 455014 480 6 mask_rev[19]
port 541 nsew signal input
rlabel metal2 s 367190 0 367246 480 6 mask_rev[1]
port 542 nsew signal input
rlabel metal2 s 459834 0 459890 480 6 mask_rev[20]
port 543 nsew signal input
rlabel metal2 s 464710 0 464766 480 6 mask_rev[21]
port 544 nsew signal input
rlabel metal2 s 469586 0 469642 480 6 mask_rev[22]
port 545 nsew signal input
rlabel metal2 s 474462 0 474518 480 6 mask_rev[23]
port 546 nsew signal input
rlabel metal2 s 479338 0 479394 480 6 mask_rev[24]
port 547 nsew signal input
rlabel metal2 s 484214 0 484270 480 6 mask_rev[25]
port 548 nsew signal input
rlabel metal2 s 489090 0 489146 480 6 mask_rev[26]
port 549 nsew signal input
rlabel metal2 s 493966 0 494022 480 6 mask_rev[27]
port 550 nsew signal input
rlabel metal2 s 498842 0 498898 480 6 mask_rev[28]
port 551 nsew signal input
rlabel metal2 s 503718 0 503774 480 6 mask_rev[29]
port 552 nsew signal input
rlabel metal2 s 372066 0 372122 480 6 mask_rev[2]
port 553 nsew signal input
rlabel metal2 s 508594 0 508650 480 6 mask_rev[30]
port 554 nsew signal input
rlabel metal2 s 513470 0 513526 480 6 mask_rev[31]
port 555 nsew signal input
rlabel metal2 s 376942 0 376998 480 6 mask_rev[3]
port 556 nsew signal input
rlabel metal2 s 381818 0 381874 480 6 mask_rev[4]
port 557 nsew signal input
rlabel metal2 s 386694 0 386750 480 6 mask_rev[5]
port 558 nsew signal input
rlabel metal2 s 391570 0 391626 480 6 mask_rev[6]
port 559 nsew signal input
rlabel metal2 s 396446 0 396502 480 6 mask_rev[7]
port 560 nsew signal input
rlabel metal2 s 401322 0 401378 480 6 mask_rev[8]
port 561 nsew signal input
rlabel metal2 s 406198 0 406254 480 6 mask_rev[9]
port 562 nsew signal input
rlabel metal3 s 0 23672 480 23792 6 por
port 563 nsew signal input
rlabel metal3 s 0 22040 480 22160 6 porb
port 564 nsew signal input
rlabel metal2 s 6366 0 6422 480 6 resetb
port 565 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 520000 320000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 219350330
string GDS_FILE /home/hosni/caravel_openframe_project/openlane/picosoc/runs/23_08_29_13_31/results/signoff/picosoc.magic.gds
string GDS_START 18154750
<< end >>

